module InHandle(
	input wire			nReset,                                                      // Common to all
	input wire			Clk,                                                        // Common to all
	output reg	[7:0]	Pixel,
	output reg			Frame,
	output reg			Line
);

	parameter COLS = 75;
	parameter ROWS = 75;
	
	reg [7:0] col;
	reg [7:0] row;
	
	always @ (posedge Clk or negedge nReset) begin
		if(!nReset) begin   
			Frame <= 0;
	    	Line  <= 0;							
			row <= ROWS-1;
			col <= COLS-1;						// Zero on first pixel	
		end else begin
			if(col == (COLS-1)) begin			// Get ready for next column
	    		Line <= 1;
				col <= 0;
				row <= row + 1;
				if(row == (ROWS-1)) begin		// Get ready for next row
					Frame <= 1;
					row <= 0;
				end
			end else begin
				Line <= 0;
				Frame <= 0;
				col = col + 1;
			end
		end
	end

	always @ (*) begin
		case(col + (row*COLS))


			0: Pixel = 161;
			1: Pixel = 159;
			2: Pixel = 156;
			3: Pixel = 154;
			4: Pixel = 154;
			5: Pixel = 160;
			6: Pixel = 170;
			7: Pixel = 170;
			8: Pixel = 145;
			9: Pixel = 100;
			10: Pixel = 96;
			11: Pixel = 106;
			12: Pixel = 106;
			13: Pixel = 107;
			14: Pixel = 106;
			15: Pixel = 110;
			16: Pixel = 119;
			17: Pixel = 124;
			18: Pixel = 128;
			19: Pixel = 131;
			20: Pixel = 131;
			21: Pixel = 129;
			22: Pixel = 130;
			23: Pixel = 132;
			24: Pixel = 133;
			25: Pixel = 134;
			26: Pixel = 132;
			27: Pixel = 132;
			28: Pixel = 134;
			29: Pixel = 134;
			30: Pixel = 134;
			31: Pixel = 131;
			32: Pixel = 130;
			33: Pixel = 132;
			34: Pixel = 130;
			35: Pixel = 133;
			36: Pixel = 132;
			37: Pixel = 134;
			38: Pixel = 130;
			39: Pixel = 129;
			40: Pixel = 129;
			41: Pixel = 129;
			42: Pixel = 129;
			43: Pixel = 127;
			44: Pixel = 125;
			45: Pixel = 119;
			46: Pixel = 106;
			47: Pixel = 121;
			48: Pixel = 149;
			49: Pixel = 159;
			50: Pixel = 153;
			51: Pixel = 152;
			52: Pixel = 154;
			53: Pixel = 154;
			54: Pixel = 152;
			55: Pixel = 152;
			56: Pixel = 155;
			57: Pixel = 157;
			58: Pixel = 154;
			59: Pixel = 194;
			60: Pixel = 223;
			61: Pixel = 191;
			62: Pixel = 104;
			63: Pixel = 115;
			64: Pixel = 121;
			65: Pixel = 121;
			66: Pixel = 121;
			67: Pixel = 121;
			68: Pixel = 124;
			69: Pixel = 123;
			70: Pixel = 123;
			71: Pixel = 126;
			72: Pixel = 119;
			73: Pixel = 129;
			74: Pixel = 145;
			75: Pixel = 157;
			76: Pixel = 156;
			77: Pixel = 155;
			78: Pixel = 154;
			79: Pixel = 153;
			80: Pixel = 162;
			81: Pixel = 170;
			82: Pixel = 167;
			83: Pixel = 139;
			84: Pixel = 97;
			85: Pixel = 92;
			86: Pixel = 103;
			87: Pixel = 105;
			88: Pixel = 104;
			89: Pixel = 103;
			90: Pixel = 110;
			91: Pixel = 119;
			92: Pixel = 124;
			93: Pixel = 126;
			94: Pixel = 128;
			95: Pixel = 129;
			96: Pixel = 131;
			97: Pixel = 129;
			98: Pixel = 131;
			99: Pixel = 132;
			100: Pixel = 133;
			101: Pixel = 131;
			102: Pixel = 132;
			103: Pixel = 131;
			104: Pixel = 131;
			105: Pixel = 131;
			106: Pixel = 130;
			107: Pixel = 128;
			108: Pixel = 130;
			109: Pixel = 129;
			110: Pixel = 132;
			111: Pixel = 130;
			112: Pixel = 130;
			113: Pixel = 130;
			114: Pixel = 128;
			115: Pixel = 127;
			116: Pixel = 127;
			117: Pixel = 128;
			118: Pixel = 127;
			119: Pixel = 125;
			120: Pixel = 119;
			121: Pixel = 108;
			122: Pixel = 110;
			123: Pixel = 139;
			124: Pixel = 156;
			125: Pixel = 157;
			126: Pixel = 154;
			127: Pixel = 157;
			128: Pixel = 156;
			129: Pixel = 154;
			130: Pixel = 154;
			131: Pixel = 153;
			132: Pixel = 154;
			133: Pixel = 150;
			134: Pixel = 171;
			135: Pixel = 215;
			136: Pixel = 217;
			137: Pixel = 137;
			138: Pixel = 104;
			139: Pixel = 119;
			140: Pixel = 120;
			141: Pixel = 120;
			142: Pixel = 121;
			143: Pixel = 122;
			144: Pixel = 123;
			145: Pixel = 123;
			146: Pixel = 125;
			147: Pixel = 133;
			148: Pixel = 98;
			149: Pixel = 53;
			150: Pixel = 156;
			151: Pixel = 156;
			152: Pixel = 157;
			153: Pixel = 154;
			154: Pixel = 158;
			155: Pixel = 167;
			156: Pixel = 166;
			157: Pixel = 161;
			158: Pixel = 138;
			159: Pixel = 98;
			160: Pixel = 92;
			161: Pixel = 104;
			162: Pixel = 106;
			163: Pixel = 104;
			164: Pixel = 102;
			165: Pixel = 110;
			166: Pixel = 117;
			167: Pixel = 123;
			168: Pixel = 126;
			169: Pixel = 128;
			170: Pixel = 130;
			171: Pixel = 131;
			172: Pixel = 130;
			173: Pixel = 130;
			174: Pixel = 132;
			175: Pixel = 133;
			176: Pixel = 132;
			177: Pixel = 131;
			178: Pixel = 131;
			179: Pixel = 132;
			180: Pixel = 132;
			181: Pixel = 132;
			182: Pixel = 130;
			183: Pixel = 130;
			184: Pixel = 129;
			185: Pixel = 134;
			186: Pixel = 134;
			187: Pixel = 130;
			188: Pixel = 131;
			189: Pixel = 129;
			190: Pixel = 128;
			191: Pixel = 127;
			192: Pixel = 128;
			193: Pixel = 128;
			194: Pixel = 127;
			195: Pixel = 120;
			196: Pixel = 114;
			197: Pixel = 104;
			198: Pixel = 125;
			199: Pixel = 152;
			200: Pixel = 160;
			201: Pixel = 160;
			202: Pixel = 161;
			203: Pixel = 161;
			204: Pixel = 157;
			205: Pixel = 156;
			206: Pixel = 154;
			207: Pixel = 152;
			208: Pixel = 151;
			209: Pixel = 148;
			210: Pixel = 192;
			211: Pixel = 224;
			212: Pixel = 197;
			213: Pixel = 109;
			214: Pixel = 112;
			215: Pixel = 119;
			216: Pixel = 121;
			217: Pixel = 121;
			218: Pixel = 123;
			219: Pixel = 124;
			220: Pixel = 127;
			221: Pixel = 136;
			222: Pixel = 94;
			223: Pixel = 45;
			224: Pixel = 45;
			225: Pixel = 155;
			226: Pixel = 157;
			227: Pixel = 158;
			228: Pixel = 155;
			229: Pixel = 163;
			230: Pixel = 166;
			231: Pixel = 161;
			232: Pixel = 160;
			233: Pixel = 141;
			234: Pixel = 98;
			235: Pixel = 91;
			236: Pixel = 104;
			237: Pixel = 105;
			238: Pixel = 103;
			239: Pixel = 103;
			240: Pixel = 109;
			241: Pixel = 117;
			242: Pixel = 122;
			243: Pixel = 125;
			244: Pixel = 128;
			245: Pixel = 129;
			246: Pixel = 129;
			247: Pixel = 129;
			248: Pixel = 130;
			249: Pixel = 130;
			250: Pixel = 131;
			251: Pixel = 130;
			252: Pixel = 130;
			253: Pixel = 132;
			254: Pixel = 129;
			255: Pixel = 128;
			256: Pixel = 128;
			257: Pixel = 129;
			258: Pixel = 127;
			259: Pixel = 127;
			260: Pixel = 130;
			261: Pixel = 133;
			262: Pixel = 130;
			263: Pixel = 130;
			264: Pixel = 128;
			265: Pixel = 127;
			266: Pixel = 126;
			267: Pixel = 127;
			268: Pixel = 127;
			269: Pixel = 126;
			270: Pixel = 123;
			271: Pixel = 115;
			272: Pixel = 105;
			273: Pixel = 117;
			274: Pixel = 147;
			275: Pixel = 160;
			276: Pixel = 162;
			277: Pixel = 160;
			278: Pixel = 160;
			279: Pixel = 158;
			280: Pixel = 156;
			281: Pixel = 154;
			282: Pixel = 152;
			283: Pixel = 152;
			284: Pixel = 146;
			285: Pixel = 159;
			286: Pixel = 211;
			287: Pixel = 225;
			288: Pixel = 156;
			289: Pixel = 101;
			290: Pixel = 119;
			291: Pixel = 122;
			292: Pixel = 121;
			293: Pixel = 122;
			294: Pixel = 127;
			295: Pixel = 138;
			296: Pixel = 94;
			297: Pixel = 42;
			298: Pixel = 46;
			299: Pixel = 51;
			300: Pixel = 157;
			301: Pixel = 158;
			302: Pixel = 159;
			303: Pixel = 162;
			304: Pixel = 168;
			305: Pixel = 164;
			306: Pixel = 157;
			307: Pixel = 161;
			308: Pixel = 140;
			309: Pixel = 95;
			310: Pixel = 91;
			311: Pixel = 103;
			312: Pixel = 106;
			313: Pixel = 103;
			314: Pixel = 103;
			315: Pixel = 108;
			316: Pixel = 117;
			317: Pixel = 122;
			318: Pixel = 125;
			319: Pixel = 127;
			320: Pixel = 127;
			321: Pixel = 127;
			322: Pixel = 129;
			323: Pixel = 129;
			324: Pixel = 130;
			325: Pixel = 130;
			326: Pixel = 129;
			327: Pixel = 129;
			328: Pixel = 133;
			329: Pixel = 128;
			330: Pixel = 122;
			331: Pixel = 122;
			332: Pixel = 126;
			333: Pixel = 126;
			334: Pixel = 125;
			335: Pixel = 127;
			336: Pixel = 129;
			337: Pixel = 131;
			338: Pixel = 129;
			339: Pixel = 126;
			340: Pixel = 127;
			341: Pixel = 126;
			342: Pixel = 126;
			343: Pixel = 126;
			344: Pixel = 127;
			345: Pixel = 122;
			346: Pixel = 115;
			347: Pixel = 107;
			348: Pixel = 119;
			349: Pixel = 142;
			350: Pixel = 157;
			351: Pixel = 160;
			352: Pixel = 158;
			353: Pixel = 158;
			354: Pixel = 157;
			355: Pixel = 156;
			356: Pixel = 155;
			357: Pixel = 155;
			358: Pixel = 154;
			359: Pixel = 151;
			360: Pixel = 142;
			361: Pixel = 183;
			362: Pixel = 222;
			363: Pixel = 212;
			364: Pixel = 122;
			365: Pixel = 111;
			366: Pixel = 122;
			367: Pixel = 121;
			368: Pixel = 122;
			369: Pixel = 135;
			370: Pixel = 91;
			371: Pixel = 40;
			372: Pixel = 47;
			373: Pixel = 49;
			374: Pixel = 53;
			375: Pixel = 159;
			376: Pixel = 160;
			377: Pixel = 164;
			378: Pixel = 167;
			379: Pixel = 166;
			380: Pixel = 161;
			381: Pixel = 158;
			382: Pixel = 161;
			383: Pixel = 139;
			384: Pixel = 94;
			385: Pixel = 90;
			386: Pixel = 103;
			387: Pixel = 103;
			388: Pixel = 102;
			389: Pixel = 102;
			390: Pixel = 108;
			391: Pixel = 116;
			392: Pixel = 120;
			393: Pixel = 122;
			394: Pixel = 125;
			395: Pixel = 127;
			396: Pixel = 125;
			397: Pixel = 126;
			398: Pixel = 129;
			399: Pixel = 128;
			400: Pixel = 128;
			401: Pixel = 130;
			402: Pixel = 129;
			403: Pixel = 129;
			404: Pixel = 126;
			405: Pixel = 123;
			406: Pixel = 121;
			407: Pixel = 120;
			408: Pixel = 118;
			409: Pixel = 116;
			410: Pixel = 123;
			411: Pixel = 129;
			412: Pixel = 132;
			413: Pixel = 129;
			414: Pixel = 127;
			415: Pixel = 128;
			416: Pixel = 126;
			417: Pixel = 125;
			418: Pixel = 126;
			419: Pixel = 126;
			420: Pixel = 121;
			421: Pixel = 117;
			422: Pixel = 109;
			423: Pixel = 117;
			424: Pixel = 138;
			425: Pixel = 151;
			426: Pixel = 156;
			427: Pixel = 157;
			428: Pixel = 157;
			429: Pixel = 156;
			430: Pixel = 155;
			431: Pixel = 156;
			432: Pixel = 156;
			433: Pixel = 154;
			434: Pixel = 152;
			435: Pixel = 144;
			436: Pixel = 150;
			437: Pixel = 208;
			438: Pixel = 229;
			439: Pixel = 180;
			440: Pixel = 101;
			441: Pixel = 115;
			442: Pixel = 121;
			443: Pixel = 134;
			444: Pixel = 90;
			445: Pixel = 38;
			446: Pixel = 50;
			447: Pixel = 55;
			448: Pixel = 51;
			449: Pixel = 48;
			450: Pixel = 161;
			451: Pixel = 161;
			452: Pixel = 167;
			453: Pixel = 160;
			454: Pixel = 155;
			455: Pixel = 159;
			456: Pixel = 160;
			457: Pixel = 161;
			458: Pixel = 139;
			459: Pixel = 92;
			460: Pixel = 89;
			461: Pixel = 103;
			462: Pixel = 103;
			463: Pixel = 103;
			464: Pixel = 102;
			465: Pixel = 108;
			466: Pixel = 117;
			467: Pixel = 120;
			468: Pixel = 123;
			469: Pixel = 124;
			470: Pixel = 125;
			471: Pixel = 125;
			472: Pixel = 128;
			473: Pixel = 127;
			474: Pixel = 127;
			475: Pixel = 129;
			476: Pixel = 129;
			477: Pixel = 127;
			478: Pixel = 127;
			479: Pixel = 127;
			480: Pixel = 129;
			481: Pixel = 128;
			482: Pixel = 138;
			483: Pixel = 140;
			484: Pixel = 137;
			485: Pixel = 128;
			486: Pixel = 120;
			487: Pixel = 119;
			488: Pixel = 125;
			489: Pixel = 127;
			490: Pixel = 129;
			491: Pixel = 127;
			492: Pixel = 126;
			493: Pixel = 126;
			494: Pixel = 125;
			495: Pixel = 120;
			496: Pixel = 116;
			497: Pixel = 110;
			498: Pixel = 115;
			499: Pixel = 136;
			500: Pixel = 146;
			501: Pixel = 151;
			502: Pixel = 155;
			503: Pixel = 155;
			504: Pixel = 154;
			505: Pixel = 153;
			506: Pixel = 154;
			507: Pixel = 154;
			508: Pixel = 150;
			509: Pixel = 146;
			510: Pixel = 145;
			511: Pixel = 137;
			512: Pixel = 178;
			513: Pixel = 223;
			514: Pixel = 222;
			515: Pixel = 133;
			516: Pixel = 101;
			517: Pixel = 126;
			518: Pixel = 91;
			519: Pixel = 40;
			520: Pixel = 46;
			521: Pixel = 57;
			522: Pixel = 55;
			523: Pixel = 47;
			524: Pixel = 45;
			525: Pixel = 159;
			526: Pixel = 164;
			527: Pixel = 165;
			528: Pixel = 145;
			529: Pixel = 143;
			530: Pixel = 161;
			531: Pixel = 162;
			532: Pixel = 162;
			533: Pixel = 141;
			534: Pixel = 93;
			535: Pixel = 88;
			536: Pixel = 101;
			537: Pixel = 104;
			538: Pixel = 103;
			539: Pixel = 104;
			540: Pixel = 111;
			541: Pixel = 118;
			542: Pixel = 121;
			543: Pixel = 124;
			544: Pixel = 126;
			545: Pixel = 126;
			546: Pixel = 128;
			547: Pixel = 129;
			548: Pixel = 128;
			549: Pixel = 125;
			550: Pixel = 128;
			551: Pixel = 128;
			552: Pixel = 128;
			553: Pixel = 140;
			554: Pixel = 144;
			555: Pixel = 147;
			556: Pixel = 161;
			557: Pixel = 173;
			558: Pixel = 182;
			559: Pixel = 180;
			560: Pixel = 178;
			561: Pixel = 170;
			562: Pixel = 146;
			563: Pixel = 120;
			564: Pixel = 117;
			565: Pixel = 129;
			566: Pixel = 129;
			567: Pixel = 126;
			568: Pixel = 125;
			569: Pixel = 124;
			570: Pixel = 120;
			571: Pixel = 115;
			572: Pixel = 109;
			573: Pixel = 113;
			574: Pixel = 137;
			575: Pixel = 144;
			576: Pixel = 145;
			577: Pixel = 151;
			578: Pixel = 154;
			579: Pixel = 151;
			580: Pixel = 152;
			581: Pixel = 152;
			582: Pixel = 148;
			583: Pixel = 145;
			584: Pixel = 142;
			585: Pixel = 141;
			586: Pixel = 140;
			587: Pixel = 146;
			588: Pixel = 202;
			589: Pixel = 229;
			590: Pixel = 195;
			591: Pixel = 120;
			592: Pixel = 88;
			593: Pixel = 39;
			594: Pixel = 46;
			595: Pixel = 52;
			596: Pixel = 55;
			597: Pixel = 50;
			598: Pixel = 46;
			599: Pixel = 46;
			600: Pixel = 162;
			601: Pixel = 169;
			602: Pixel = 154;
			603: Pixel = 123;
			604: Pixel = 139;
			605: Pixel = 164;
			606: Pixel = 164;
			607: Pixel = 164;
			608: Pixel = 141;
			609: Pixel = 90;
			610: Pixel = 85;
			611: Pixel = 98;
			612: Pixel = 100;
			613: Pixel = 101;
			614: Pixel = 104;
			615: Pixel = 110;
			616: Pixel = 117;
			617: Pixel = 121;
			618: Pixel = 123;
			619: Pixel = 123;
			620: Pixel = 124;
			621: Pixel = 127;
			622: Pixel = 126;
			623: Pixel = 127;
			624: Pixel = 134;
			625: Pixel = 137;
			626: Pixel = 126;
			627: Pixel = 134;
			628: Pixel = 142;
			629: Pixel = 144;
			630: Pixel = 149;
			631: Pixel = 157;
			632: Pixel = 165;
			633: Pixel = 172;
			634: Pixel = 174;
			635: Pixel = 179;
			636: Pixel = 189;
			637: Pixel = 198;
			638: Pixel = 184;
			639: Pixel = 136;
			640: Pixel = 113;
			641: Pixel = 123;
			642: Pixel = 125;
			643: Pixel = 123;
			644: Pixel = 120;
			645: Pixel = 115;
			646: Pixel = 112;
			647: Pixel = 106;
			648: Pixel = 113;
			649: Pixel = 138;
			650: Pixel = 146;
			651: Pixel = 144;
			652: Pixel = 148;
			653: Pixel = 151;
			654: Pixel = 151;
			655: Pixel = 146;
			656: Pixel = 145;
			657: Pixel = 145;
			658: Pixel = 143;
			659: Pixel = 140;
			660: Pixel = 139;
			661: Pixel = 141;
			662: Pixel = 135;
			663: Pixel = 163;
			664: Pixel = 219;
			665: Pixel = 238;
			666: Pixel = 145;
			667: Pixel = 32;
			668: Pixel = 46;
			669: Pixel = 52;
			670: Pixel = 54;
			671: Pixel = 49;
			672: Pixel = 50;
			673: Pixel = 48;
			674: Pixel = 47;
			675: Pixel = 170;
			676: Pixel = 166;
			677: Pixel = 131;
			678: Pixel = 95;
			679: Pixel = 142;
			680: Pixel = 166;
			681: Pixel = 164;
			682: Pixel = 163;
			683: Pixel = 142;
			684: Pixel = 89;
			685: Pixel = 80;
			686: Pixel = 94;
			687: Pixel = 97;
			688: Pixel = 99;
			689: Pixel = 102;
			690: Pixel = 106;
			691: Pixel = 113;
			692: Pixel = 117;
			693: Pixel = 120;
			694: Pixel = 122;
			695: Pixel = 124;
			696: Pixel = 123;
			697: Pixel = 127;
			698: Pixel = 129;
			699: Pixel = 128;
			700: Pixel = 126;
			701: Pixel = 121;
			702: Pixel = 130;
			703: Pixel = 129;
			704: Pixel = 135;
			705: Pixel = 142;
			706: Pixel = 151;
			707: Pixel = 161;
			708: Pixel = 170;
			709: Pixel = 179;
			710: Pixel = 184;
			711: Pixel = 185;
			712: Pixel = 187;
			713: Pixel = 197;
			714: Pixel = 200;
			715: Pixel = 160;
			716: Pixel = 112;
			717: Pixel = 111;
			718: Pixel = 119;
			719: Pixel = 118;
			720: Pixel = 114;
			721: Pixel = 110;
			722: Pixel = 103;
			723: Pixel = 111;
			724: Pixel = 138;
			725: Pixel = 148;
			726: Pixel = 144;
			727: Pixel = 145;
			728: Pixel = 145;
			729: Pixel = 150;
			730: Pixel = 145;
			731: Pixel = 140;
			732: Pixel = 144;
			733: Pixel = 143;
			734: Pixel = 142;
			735: Pixel = 140;
			736: Pixel = 142;
			737: Pixel = 143;
			738: Pixel = 138;
			739: Pixel = 197;
			740: Pixel = 228;
			741: Pixel = 81;
			742: Pixel = 34;
			743: Pixel = 51;
			744: Pixel = 55;
			745: Pixel = 49;
			746: Pixel = 47;
			747: Pixel = 48;
			748: Pixel = 48;
			749: Pixel = 47;
			750: Pixel = 171;
			751: Pixel = 154;
			752: Pixel = 97;
			753: Pixel = 86;
			754: Pixel = 142;
			755: Pixel = 166;
			756: Pixel = 165;
			757: Pixel = 161;
			758: Pixel = 138;
			759: Pixel = 86;
			760: Pixel = 79;
			761: Pixel = 96;
			762: Pixel = 100;
			763: Pixel = 100;
			764: Pixel = 100;
			765: Pixel = 105;
			766: Pixel = 112;
			767: Pixel = 114;
			768: Pixel = 118;
			769: Pixel = 120;
			770: Pixel = 123;
			771: Pixel = 123;
			772: Pixel = 131;
			773: Pixel = 114;
			774: Pixel = 112;
			775: Pixel = 119;
			776: Pixel = 124;
			777: Pixel = 129;
			778: Pixel = 132;
			779: Pixel = 134;
			780: Pixel = 135;
			781: Pixel = 143;
			782: Pixel = 157;
			783: Pixel = 170;
			784: Pixel = 176;
			785: Pixel = 182;
			786: Pixel = 188;
			787: Pixel = 191;
			788: Pixel = 195;
			789: Pixel = 194;
			790: Pixel = 202;
			791: Pixel = 182;
			792: Pixel = 115;
			793: Pixel = 97;
			794: Pixel = 113;
			795: Pixel = 111;
			796: Pixel = 108;
			797: Pixel = 103;
			798: Pixel = 109;
			799: Pixel = 141;
			800: Pixel = 153;
			801: Pixel = 150;
			802: Pixel = 141;
			803: Pixel = 134;
			804: Pixel = 140;
			805: Pixel = 148;
			806: Pixel = 142;
			807: Pixel = 145;
			808: Pixel = 143;
			809: Pixel = 141;
			810: Pixel = 143;
			811: Pixel = 144;
			812: Pixel = 145;
			813: Pixel = 146;
			814: Pixel = 166;
			815: Pixel = 94;
			816: Pixel = 33;
			817: Pixel = 49;
			818: Pixel = 52;
			819: Pixel = 49;
			820: Pixel = 50;
			821: Pixel = 51;
			822: Pixel = 50;
			823: Pixel = 54;
			824: Pixel = 43;
			825: Pixel = 163;
			826: Pixel = 128;
			827: Pixel = 79;
			828: Pixel = 94;
			829: Pixel = 142;
			830: Pixel = 166;
			831: Pixel = 167;
			832: Pixel = 162;
			833: Pixel = 138;
			834: Pixel = 85;
			835: Pixel = 80;
			836: Pixel = 97;
			837: Pixel = 99;
			838: Pixel = 99;
			839: Pixel = 100;
			840: Pixel = 105;
			841: Pixel = 112;
			842: Pixel = 115;
			843: Pixel = 118;
			844: Pixel = 121;
			845: Pixel = 120;
			846: Pixel = 128;
			847: Pixel = 126;
			848: Pixel = 107;
			849: Pixel = 114;
			850: Pixel = 118;
			851: Pixel = 124;
			852: Pixel = 126;
			853: Pixel = 130;
			854: Pixel = 135;
			855: Pixel = 135;
			856: Pixel = 141;
			857: Pixel = 149;
			858: Pixel = 164;
			859: Pixel = 181;
			860: Pixel = 185;
			861: Pixel = 189;
			862: Pixel = 191;
			863: Pixel = 190;
			864: Pixel = 192;
			865: Pixel = 197;
			866: Pixel = 211;
			867: Pixel = 222;
			868: Pixel = 153;
			869: Pixel = 87;
			870: Pixel = 108;
			871: Pixel = 103;
			872: Pixel = 100;
			873: Pixel = 108;
			874: Pixel = 142;
			875: Pixel = 155;
			876: Pixel = 154;
			877: Pixel = 145;
			878: Pixel = 113;
			879: Pixel = 115;
			880: Pixel = 145;
			881: Pixel = 146;
			882: Pixel = 145;
			883: Pixel = 144;
			884: Pixel = 143;
			885: Pixel = 144;
			886: Pixel = 145;
			887: Pixel = 146;
			888: Pixel = 160;
			889: Pixel = 95;
			890: Pixel = 32;
			891: Pixel = 46;
			892: Pixel = 52;
			893: Pixel = 50;
			894: Pixel = 47;
			895: Pixel = 52;
			896: Pixel = 48;
			897: Pixel = 64;
			898: Pixel = 49;
			899: Pixel = 122;
			900: Pixel = 145;
			901: Pixel = 96;
			902: Pixel = 82;
			903: Pixel = 96;
			904: Pixel = 141;
			905: Pixel = 165;
			906: Pixel = 167;
			907: Pixel = 162;
			908: Pixel = 136;
			909: Pixel = 87;
			910: Pixel = 82;
			911: Pixel = 96;
			912: Pixel = 99;
			913: Pixel = 101;
			914: Pixel = 101;
			915: Pixel = 105;
			916: Pixel = 112;
			917: Pixel = 115;
			918: Pixel = 119;
			919: Pixel = 121;
			920: Pixel = 123;
			921: Pixel = 122;
			922: Pixel = 107;
			923: Pixel = 112;
			924: Pixel = 119;
			925: Pixel = 120;
			926: Pixel = 118;
			927: Pixel = 122;
			928: Pixel = 130;
			929: Pixel = 135;
			930: Pixel = 134;
			931: Pixel = 139;
			932: Pixel = 148;
			933: Pixel = 164;
			934: Pixel = 182;
			935: Pixel = 186;
			936: Pixel = 179;
			937: Pixel = 185;
			938: Pixel = 198;
			939: Pixel = 207;
			940: Pixel = 210;
			941: Pixel = 207;
			942: Pixel = 214;
			943: Pixel = 226;
			944: Pixel = 117;
			945: Pixel = 84;
			946: Pixel = 103;
			947: Pixel = 96;
			948: Pixel = 106;
			949: Pixel = 140;
			950: Pixel = 154;
			951: Pixel = 153;
			952: Pixel = 150;
			953: Pixel = 104;
			954: Pixel = 70;
			955: Pixel = 126;
			956: Pixel = 148;
			957: Pixel = 144;
			958: Pixel = 144;
			959: Pixel = 143;
			960: Pixel = 144;
			961: Pixel = 142;
			962: Pixel = 155;
			963: Pixel = 124;
			964: Pixel = 39;
			965: Pixel = 44;
			966: Pixel = 54;
			967: Pixel = 52;
			968: Pixel = 46;
			969: Pixel = 51;
			970: Pixel = 48;
			971: Pixel = 61;
			972: Pixel = 67;
			973: Pixel = 113;
			974: Pixel = 156;
			975: Pixel = 110;
			976: Pixel = 86;
			977: Pixel = 88;
			978: Pixel = 94;
			979: Pixel = 140;
			980: Pixel = 164;
			981: Pixel = 166;
			982: Pixel = 162;
			983: Pixel = 136;
			984: Pixel = 87;
			985: Pixel = 83;
			986: Pixel = 97;
			987: Pixel = 99;
			988: Pixel = 101;
			989: Pixel = 100;
			990: Pixel = 105;
			991: Pixel = 112;
			992: Pixel = 116;
			993: Pixel = 119;
			994: Pixel = 121;
			995: Pixel = 123;
			996: Pixel = 109;
			997: Pixel = 110;
			998: Pixel = 116;
			999: Pixel = 117;
			1000: Pixel = 113;
			1001: Pixel = 119;
			1002: Pixel = 127;
			1003: Pixel = 134;
			1004: Pixel = 139;
			1005: Pixel = 143;
			1006: Pixel = 142;
			1007: Pixel = 145;
			1008: Pixel = 164;
			1009: Pixel = 171;
			1010: Pixel = 169;
			1011: Pixel = 188;
			1012: Pixel = 204;
			1013: Pixel = 209;
			1014: Pixel = 203;
			1015: Pixel = 202;
			1016: Pixel = 205;
			1017: Pixel = 207;
			1018: Pixel = 220;
			1019: Pixel = 210;
			1020: Pixel = 88;
			1021: Pixel = 79;
			1022: Pixel = 93;
			1023: Pixel = 104;
			1024: Pixel = 140;
			1025: Pixel = 155;
			1026: Pixel = 153;
			1027: Pixel = 151;
			1028: Pixel = 112;
			1029: Pixel = 45;
			1030: Pixel = 94;
			1031: Pixel = 142;
			1032: Pixel = 147;
			1033: Pixel = 143;
			1034: Pixel = 143;
			1035: Pixel = 143;
			1036: Pixel = 148;
			1037: Pixel = 147;
			1038: Pixel = 57;
			1039: Pixel = 44;
			1040: Pixel = 52;
			1041: Pixel = 54;
			1042: Pixel = 47;
			1043: Pixel = 53;
			1044: Pixel = 49;
			1045: Pixel = 53;
			1046: Pixel = 71;
			1047: Pixel = 113;
			1048: Pixel = 150;
			1049: Pixel = 144;
			1050: Pixel = 87;
			1051: Pixel = 90;
			1052: Pixel = 89;
			1053: Pixel = 93;
			1054: Pixel = 138;
			1055: Pixel = 162;
			1056: Pixel = 166;
			1057: Pixel = 162;
			1058: Pixel = 136;
			1059: Pixel = 88;
			1060: Pixel = 81;
			1061: Pixel = 98;
			1062: Pixel = 99;
			1063: Pixel = 99;
			1064: Pixel = 101;
			1065: Pixel = 104;
			1066: Pixel = 112;
			1067: Pixel = 117;
			1068: Pixel = 118;
			1069: Pixel = 124;
			1070: Pixel = 117;
			1071: Pixel = 111;
			1072: Pixel = 113;
			1073: Pixel = 115;
			1074: Pixel = 116;
			1075: Pixel = 118;
			1076: Pixel = 126;
			1077: Pixel = 131;
			1078: Pixel = 137;
			1079: Pixel = 139;
			1080: Pixel = 141;
			1081: Pixel = 138;
			1082: Pixel = 143;
			1083: Pixel = 153;
			1084: Pixel = 164;
			1085: Pixel = 192;
			1086: Pixel = 205;
			1087: Pixel = 202;
			1088: Pixel = 199;
			1089: Pixel = 197;
			1090: Pixel = 201;
			1091: Pixel = 203;
			1092: Pixel = 206;
			1093: Pixel = 207;
			1094: Pixel = 218;
			1095: Pixel = 203;
			1096: Pixel = 104;
			1097: Pixel = 71;
			1098: Pixel = 103;
			1099: Pixel = 141;
			1100: Pixel = 155;
			1101: Pixel = 153;
			1102: Pixel = 153;
			1103: Pixel = 112;
			1104: Pixel = 45;
			1105: Pixel = 60;
			1106: Pixel = 120;
			1107: Pixel = 149;
			1108: Pixel = 145;
			1109: Pixel = 142;
			1110: Pixel = 145;
			1111: Pixel = 158;
			1112: Pixel = 88;
			1113: Pixel = 32;
			1114: Pixel = 51;
			1115: Pixel = 57;
			1116: Pixel = 47;
			1117: Pixel = 50;
			1118: Pixel = 51;
			1119: Pixel = 52;
			1120: Pixel = 54;
			1121: Pixel = 103;
			1122: Pixel = 149;
			1123: Pixel = 147;
			1124: Pixel = 162;
			1125: Pixel = 89;
			1126: Pixel = 93;
			1127: Pixel = 90;
			1128: Pixel = 96;
			1129: Pixel = 138;
			1130: Pixel = 161;
			1131: Pixel = 165;
			1132: Pixel = 162;
			1133: Pixel = 137;
			1134: Pixel = 88;
			1135: Pixel = 80;
			1136: Pixel = 95;
			1137: Pixel = 99;
			1138: Pixel = 101;
			1139: Pixel = 100;
			1140: Pixel = 104;
			1141: Pixel = 112;
			1142: Pixel = 116;
			1143: Pixel = 118;
			1144: Pixel = 133;
			1145: Pixel = 103;
			1146: Pixel = 110;
			1147: Pixel = 113;
			1148: Pixel = 113;
			1149: Pixel = 116;
			1150: Pixel = 123;
			1151: Pixel = 133;
			1152: Pixel = 139;
			1153: Pixel = 137;
			1154: Pixel = 141;
			1155: Pixel = 135;
			1156: Pixel = 126;
			1157: Pixel = 136;
			1158: Pixel = 168;
			1159: Pixel = 195;
			1160: Pixel = 196;
			1161: Pixel = 189;
			1162: Pixel = 191;
			1163: Pixel = 198;
			1164: Pixel = 203;
			1165: Pixel = 204;
			1166: Pixel = 206;
			1167: Pixel = 207;
			1168: Pixel = 207;
			1169: Pixel = 205;
			1170: Pixel = 223;
			1171: Pixel = 208;
			1172: Pixel = 76;
			1173: Pixel = 92;
			1174: Pixel = 139;
			1175: Pixel = 154;
			1176: Pixel = 154;
			1177: Pixel = 152;
			1178: Pixel = 113;
			1179: Pixel = 51;
			1180: Pixel = 38;
			1181: Pixel = 79;
			1182: Pixel = 127;
			1183: Pixel = 140;
			1184: Pixel = 133;
			1185: Pixel = 149;
			1186: Pixel = 124;
			1187: Pixel = 39;
			1188: Pixel = 46;
			1189: Pixel = 54;
			1190: Pixel = 53;
			1191: Pixel = 50;
			1192: Pixel = 51;
			1193: Pixel = 52;
			1194: Pixel = 45;
			1195: Pixel = 86;
			1196: Pixel = 146;
			1197: Pixel = 140;
			1198: Pixel = 160;
			1199: Pixel = 165;
			1200: Pixel = 91;
			1201: Pixel = 91;
			1202: Pixel = 87;
			1203: Pixel = 92;
			1204: Pixel = 138;
			1205: Pixel = 162;
			1206: Pixel = 163;
			1207: Pixel = 163;
			1208: Pixel = 139;
			1209: Pixel = 89;
			1210: Pixel = 80;
			1211: Pixel = 94;
			1212: Pixel = 97;
			1213: Pixel = 100;
			1214: Pixel = 101;
			1215: Pixel = 107;
			1216: Pixel = 112;
			1217: Pixel = 108;
			1218: Pixel = 132;
			1219: Pixel = 142;
			1220: Pixel = 97;
			1221: Pixel = 110;
			1222: Pixel = 112;
			1223: Pixel = 115;
			1224: Pixel = 121;
			1225: Pixel = 128;
			1226: Pixel = 137;
			1227: Pixel = 134;
			1228: Pixel = 135;
			1229: Pixel = 135;
			1230: Pixel = 118;
			1231: Pixel = 134;
			1232: Pixel = 179;
			1233: Pixel = 190;
			1234: Pixel = 186;
			1235: Pixel = 183;
			1236: Pixel = 189;
			1237: Pixel = 195;
			1238: Pixel = 197;
			1239: Pixel = 204;
			1240: Pixel = 202;
			1241: Pixel = 202;
			1242: Pixel = 202;
			1243: Pixel = 204;
			1244: Pixel = 207;
			1245: Pixel = 206;
			1246: Pixel = 231;
			1247: Pixel = 160;
			1248: Pixel = 73;
			1249: Pixel = 140;
			1250: Pixel = 152;
			1251: Pixel = 153;
			1252: Pixel = 152;
			1253: Pixel = 114;
			1254: Pixel = 55;
			1255: Pixel = 42;
			1256: Pixel = 30;
			1257: Pixel = 125;
			1258: Pixel = 189;
			1259: Pixel = 182;
			1260: Pixel = 165;
			1261: Pixel = 56;
			1262: Pixel = 42;
			1263: Pixel = 54;
			1264: Pixel = 55;
			1265: Pixel = 54;
			1266: Pixel = 51;
			1267: Pixel = 52;
			1268: Pixel = 46;
			1269: Pixel = 62;
			1270: Pixel = 142;
			1271: Pixel = 142;
			1272: Pixel = 154;
			1273: Pixel = 161;
			1274: Pixel = 159;
			1275: Pixel = 89;
			1276: Pixel = 90;
			1277: Pixel = 88;
			1278: Pixel = 90;
			1279: Pixel = 136;
			1280: Pixel = 162;
			1281: Pixel = 164;
			1282: Pixel = 162;
			1283: Pixel = 138;
			1284: Pixel = 85;
			1285: Pixel = 75;
			1286: Pixel = 91;
			1287: Pixel = 96;
			1288: Pixel = 97;
			1289: Pixel = 99;
			1290: Pixel = 104;
			1291: Pixel = 110;
			1292: Pixel = 101;
			1293: Pixel = 160;
			1294: Pixel = 134;
			1295: Pixel = 96;
			1296: Pixel = 112;
			1297: Pixel = 114;
			1298: Pixel = 115;
			1299: Pixel = 124;
			1300: Pixel = 131;
			1301: Pixel = 128;
			1302: Pixel = 133;
			1303: Pixel = 130;
			1304: Pixel = 112;
			1305: Pixel = 147;
			1306: Pixel = 179;
			1307: Pixel = 180;
			1308: Pixel = 175;
			1309: Pixel = 179;
			1310: Pixel = 184;
			1311: Pixel = 190;
			1312: Pixel = 196;
			1313: Pixel = 195;
			1314: Pixel = 193;
			1315: Pixel = 197;
			1316: Pixel = 201;
			1317: Pixel = 203;
			1318: Pixel = 201;
			1319: Pixel = 206;
			1320: Pixel = 205;
			1321: Pixel = 212;
			1322: Pixel = 216;
			1323: Pixel = 94;
			1324: Pixel = 128;
			1325: Pixel = 155;
			1326: Pixel = 153;
			1327: Pixel = 153;
			1328: Pixel = 116;
			1329: Pixel = 44;
			1330: Pixel = 33;
			1331: Pixel = 126;
			1332: Pixel = 203;
			1333: Pixel = 212;
			1334: Pixel = 227;
			1335: Pixel = 220;
			1336: Pixel = 63;
			1337: Pixel = 42;
			1338: Pixel = 56;
			1339: Pixel = 53;
			1340: Pixel = 51;
			1341: Pixel = 50;
			1342: Pixel = 54;
			1343: Pixel = 47;
			1344: Pixel = 126;
			1345: Pixel = 148;
			1346: Pixel = 151;
			1347: Pixel = 163;
			1348: Pixel = 158;
			1349: Pixel = 157;
			1350: Pixel = 92;
			1351: Pixel = 94;
			1352: Pixel = 94;
			1353: Pixel = 95;
			1354: Pixel = 134;
			1355: Pixel = 163;
			1356: Pixel = 167;
			1357: Pixel = 163;
			1358: Pixel = 138;
			1359: Pixel = 85;
			1360: Pixel = 76;
			1361: Pixel = 94;
			1362: Pixel = 99;
			1363: Pixel = 100;
			1364: Pixel = 101;
			1365: Pixel = 104;
			1366: Pixel = 111;
			1367: Pixel = 108;
			1368: Pixel = 180;
			1369: Pixel = 121;
			1370: Pixel = 98;
			1371: Pixel = 108;
			1372: Pixel = 111;
			1373: Pixel = 122;
			1374: Pixel = 125;
			1375: Pixel = 120;
			1376: Pixel = 129;
			1377: Pixel = 126;
			1378: Pixel = 114;
			1379: Pixel = 154;
			1380: Pixel = 178;
			1381: Pixel = 166;
			1382: Pixel = 170;
			1383: Pixel = 178;
			1384: Pixel = 179;
			1385: Pixel = 187;
			1386: Pixel = 189;
			1387: Pixel = 185;
			1388: Pixel = 187;
			1389: Pixel = 195;
			1390: Pixel = 197;
			1391: Pixel = 196;
			1392: Pixel = 200;
			1393: Pixel = 201;
			1394: Pixel = 202;
			1395: Pixel = 204;
			1396: Pixel = 203;
			1397: Pixel = 220;
			1398: Pixel = 171;
			1399: Pixel = 118;
			1400: Pixel = 156;
			1401: Pixel = 157;
			1402: Pixel = 151;
			1403: Pixel = 91;
			1404: Pixel = 53;
			1405: Pixel = 156;
			1406: Pixel = 202;
			1407: Pixel = 206;
			1408: Pixel = 212;
			1409: Pixel = 205;
			1410: Pixel = 232;
			1411: Pixel = 100;
			1412: Pixel = 36;
			1413: Pixel = 55;
			1414: Pixel = 47;
			1415: Pixel = 45;
			1416: Pixel = 52;
			1417: Pixel = 44;
			1418: Pixel = 97;
			1419: Pixel = 154;
			1420: Pixel = 147;
			1421: Pixel = 160;
			1422: Pixel = 158;
			1423: Pixel = 157;
			1424: Pixel = 157;
			1425: Pixel = 97;
			1426: Pixel = 100;
			1427: Pixel = 97;
			1428: Pixel = 98;
			1429: Pixel = 135;
			1430: Pixel = 163;
			1431: Pixel = 167;
			1432: Pixel = 166;
			1433: Pixel = 141;
			1434: Pixel = 88;
			1435: Pixel = 81;
			1436: Pixel = 96;
			1437: Pixel = 101;
			1438: Pixel = 102;
			1439: Pixel = 101;
			1440: Pixel = 107;
			1441: Pixel = 110;
			1442: Pixel = 117;
			1443: Pixel = 184;
			1444: Pixel = 110;
			1445: Pixel = 98;
			1446: Pixel = 106;
			1447: Pixel = 113;
			1448: Pixel = 119;
			1449: Pixel = 120;
			1450: Pixel = 127;
			1451: Pixel = 126;
			1452: Pixel = 117;
			1453: Pixel = 150;
			1454: Pixel = 161;
			1455: Pixel = 156;
			1456: Pixel = 166;
			1457: Pixel = 178;
			1458: Pixel = 180;
			1459: Pixel = 180;
			1460: Pixel = 183;
			1461: Pixel = 176;
			1462: Pixel = 178;
			1463: Pixel = 187;
			1464: Pixel = 193;
			1465: Pixel = 194;
			1466: Pixel = 198;
			1467: Pixel = 198;
			1468: Pixel = 183;
			1469: Pixel = 195;
			1470: Pixel = 201;
			1471: Pixel = 202;
			1472: Pixel = 200;
			1473: Pixel = 213;
			1474: Pixel = 178;
			1475: Pixel = 147;
			1476: Pixel = 151;
			1477: Pixel = 137;
			1478: Pixel = 133;
			1479: Pixel = 186;
			1480: Pixel = 205;
			1481: Pixel = 205;
			1482: Pixel = 208;
			1483: Pixel = 200;
			1484: Pixel = 207;
			1485: Pixel = 229;
			1486: Pixel = 92;
			1487: Pixel = 39;
			1488: Pixel = 55;
			1489: Pixel = 46;
			1490: Pixel = 50;
			1491: Pixel = 45;
			1492: Pixel = 54;
			1493: Pixel = 146;
			1494: Pixel = 149;
			1495: Pixel = 159;
			1496: Pixel = 158;
			1497: Pixel = 156;
			1498: Pixel = 155;
			1499: Pixel = 155;
			1500: Pixel = 100;
			1501: Pixel = 100;
			1502: Pixel = 98;
			1503: Pixel = 101;
			1504: Pixel = 137;
			1505: Pixel = 162;
			1506: Pixel = 169;
			1507: Pixel = 170;
			1508: Pixel = 143;
			1509: Pixel = 88;
			1510: Pixel = 82;
			1511: Pixel = 97;
			1512: Pixel = 100;
			1513: Pixel = 101;
			1514: Pixel = 99;
			1515: Pixel = 106;
			1516: Pixel = 102;
			1517: Pixel = 126;
			1518: Pixel = 180;
			1519: Pixel = 111;
			1520: Pixel = 102;
			1521: Pixel = 104;
			1522: Pixel = 106;
			1523: Pixel = 114;
			1524: Pixel = 122;
			1525: Pixel = 119;
			1526: Pixel = 119;
			1527: Pixel = 146;
			1528: Pixel = 154;
			1529: Pixel = 142;
			1530: Pixel = 154;
			1531: Pixel = 171;
			1532: Pixel = 172;
			1533: Pixel = 170;
			1534: Pixel = 177;
			1535: Pixel = 170;
			1536: Pixel = 174;
			1537: Pixel = 181;
			1538: Pixel = 180;
			1539: Pixel = 181;
			1540: Pixel = 187;
			1541: Pixel = 190;
			1542: Pixel = 183;
			1543: Pixel = 181;
			1544: Pixel = 193;
			1545: Pixel = 198;
			1546: Pixel = 195;
			1547: Pixel = 194;
			1548: Pixel = 193;
			1549: Pixel = 202;
			1550: Pixel = 157;
			1551: Pixel = 156;
			1552: Pixel = 185;
			1553: Pixel = 202;
			1554: Pixel = 201;
			1555: Pixel = 204;
			1556: Pixel = 202;
			1557: Pixel = 201;
			1558: Pixel = 204;
			1559: Pixel = 215;
			1560: Pixel = 219;
			1561: Pixel = 71;
			1562: Pixel = 45;
			1563: Pixel = 51;
			1564: Pixel = 45;
			1565: Pixel = 51;
			1566: Pixel = 49;
			1567: Pixel = 114;
			1568: Pixel = 154;
			1569: Pixel = 153;
			1570: Pixel = 160;
			1571: Pixel = 157;
			1572: Pixel = 156;
			1573: Pixel = 155;
			1574: Pixel = 153;
			1575: Pixel = 100;
			1576: Pixel = 99;
			1577: Pixel = 98;
			1578: Pixel = 103;
			1579: Pixel = 138;
			1580: Pixel = 165;
			1581: Pixel = 172;
			1582: Pixel = 173;
			1583: Pixel = 145;
			1584: Pixel = 88;
			1585: Pixel = 81;
			1586: Pixel = 95;
			1587: Pixel = 99;
			1588: Pixel = 98;
			1589: Pixel = 98;
			1590: Pixel = 105;
			1591: Pixel = 94;
			1592: Pixel = 142;
			1593: Pixel = 187;
			1594: Pixel = 121;
			1595: Pixel = 106;
			1596: Pixel = 105;
			1597: Pixel = 110;
			1598: Pixel = 117;
			1599: Pixel = 120;
			1600: Pixel = 120;
			1601: Pixel = 146;
			1602: Pixel = 147;
			1603: Pixel = 136;
			1604: Pixel = 145;
			1605: Pixel = 159;
			1606: Pixel = 160;
			1607: Pixel = 171;
			1608: Pixel = 169;
			1609: Pixel = 164;
			1610: Pixel = 172;
			1611: Pixel = 175;
			1612: Pixel = 175;
			1613: Pixel = 173;
			1614: Pixel = 183;
			1615: Pixel = 183;
			1616: Pixel = 177;
			1617: Pixel = 184;
			1618: Pixel = 188;
			1619: Pixel = 190;
			1620: Pixel = 184;
			1621: Pixel = 184;
			1622: Pixel = 187;
			1623: Pixel = 177;
			1624: Pixel = 184;
			1625: Pixel = 186;
			1626: Pixel = 195;
			1627: Pixel = 201;
			1628: Pixel = 200;
			1629: Pixel = 203;
			1630: Pixel = 198;
			1631: Pixel = 201;
			1632: Pixel = 204;
			1633: Pixel = 198;
			1634: Pixel = 220;
			1635: Pixel = 200;
			1636: Pixel = 47;
			1637: Pixel = 49;
			1638: Pixel = 50;
			1639: Pixel = 47;
			1640: Pixel = 49;
			1641: Pixel = 89;
			1642: Pixel = 149;
			1643: Pixel = 149;
			1644: Pixel = 160;
			1645: Pixel = 159;
			1646: Pixel = 157;
			1647: Pixel = 157;
			1648: Pixel = 154;
			1649: Pixel = 155;
			1650: Pixel = 98;
			1651: Pixel = 98;
			1652: Pixel = 97;
			1653: Pixel = 101;
			1654: Pixel = 136;
			1655: Pixel = 167;
			1656: Pixel = 173;
			1657: Pixel = 172;
			1658: Pixel = 145;
			1659: Pixel = 89;
			1660: Pixel = 81;
			1661: Pixel = 96;
			1662: Pixel = 99;
			1663: Pixel = 99;
			1664: Pixel = 98;
			1665: Pixel = 104;
			1666: Pixel = 92;
			1667: Pixel = 152;
			1668: Pixel = 187;
			1669: Pixel = 139;
			1670: Pixel = 122;
			1671: Pixel = 104;
			1672: Pixel = 108;
			1673: Pixel = 114;
			1674: Pixel = 118;
			1675: Pixel = 140;
			1676: Pixel = 144;
			1677: Pixel = 132;
			1678: Pixel = 144;
			1679: Pixel = 152;
			1680: Pixel = 143;
			1681: Pixel = 158;
			1682: Pixel = 164;
			1683: Pixel = 164;
			1684: Pixel = 171;
			1685: Pixel = 169;
			1686: Pixel = 174;
			1687: Pixel = 171;
			1688: Pixel = 168;
			1689: Pixel = 171;
			1690: Pixel = 176;
			1691: Pixel = 180;
			1692: Pixel = 183;
			1693: Pixel = 186;
			1694: Pixel = 180;
			1695: Pixel = 179;
			1696: Pixel = 174;
			1697: Pixel = 171;
			1698: Pixel = 175;
			1699: Pixel = 187;
			1700: Pixel = 193;
			1701: Pixel = 201;
			1702: Pixel = 202;
			1703: Pixel = 198;
			1704: Pixel = 198;
			1705: Pixel = 199;
			1706: Pixel = 207;
			1707: Pixel = 181;
			1708: Pixel = 174;
			1709: Pixel = 214;
			1710: Pixel = 150;
			1711: Pixel = 33;
			1712: Pixel = 52;
			1713: Pixel = 48;
			1714: Pixel = 48;
			1715: Pixel = 53;
			1716: Pixel = 130;
			1717: Pixel = 151;
			1718: Pixel = 156;
			1719: Pixel = 161;
			1720: Pixel = 159;
			1721: Pixel = 157;
			1722: Pixel = 157;
			1723: Pixel = 157;
			1724: Pixel = 157;
			1725: Pixel = 96;
			1726: Pixel = 95;
			1727: Pixel = 95;
			1728: Pixel = 100;
			1729: Pixel = 139;
			1730: Pixel = 167;
			1731: Pixel = 171;
			1732: Pixel = 170;
			1733: Pixel = 146;
			1734: Pixel = 90;
			1735: Pixel = 83;
			1736: Pixel = 98;
			1737: Pixel = 99;
			1738: Pixel = 98;
			1739: Pixel = 98;
			1740: Pixel = 103;
			1741: Pixel = 89;
			1742: Pixel = 151;
			1743: Pixel = 185;
			1744: Pixel = 148;
			1745: Pixel = 134;
			1746: Pixel = 105;
			1747: Pixel = 102;
			1748: Pixel = 116;
			1749: Pixel = 136;
			1750: Pixel = 138;
			1751: Pixel = 127;
			1752: Pixel = 137;
			1753: Pixel = 148;
			1754: Pixel = 142;
			1755: Pixel = 150;
			1756: Pixel = 147;
			1757: Pixel = 156;
			1758: Pixel = 166;
			1759: Pixel = 166;
			1760: Pixel = 167;
			1761: Pixel = 168;
			1762: Pixel = 162;
			1763: Pixel = 161;
			1764: Pixel = 162;
			1765: Pixel = 168;
			1766: Pixel = 171;
			1767: Pixel = 176;
			1768: Pixel = 174;
			1769: Pixel = 169;
			1770: Pixel = 170;
			1771: Pixel = 167;
			1772: Pixel = 179;
			1773: Pixel = 192;
			1774: Pixel = 200;
			1775: Pixel = 199;
			1776: Pixel = 193;
			1777: Pixel = 193;
			1778: Pixel = 199;
			1779: Pixel = 200;
			1780: Pixel = 206;
			1781: Pixel = 195;
			1782: Pixel = 164;
			1783: Pixel = 154;
			1784: Pixel = 188;
			1785: Pixel = 88;
			1786: Pixel = 39;
			1787: Pixel = 52;
			1788: Pixel = 45;
			1789: Pixel = 47;
			1790: Pixel = 103;
			1791: Pixel = 151;
			1792: Pixel = 150;
			1793: Pixel = 161;
			1794: Pixel = 159;
			1795: Pixel = 158;
			1796: Pixel = 158;
			1797: Pixel = 156;
			1798: Pixel = 158;
			1799: Pixel = 156;
			1800: Pixel = 96;
			1801: Pixel = 95;
			1802: Pixel = 94;
			1803: Pixel = 103;
			1804: Pixel = 140;
			1805: Pixel = 167;
			1806: Pixel = 171;
			1807: Pixel = 171;
			1808: Pixel = 148;
			1809: Pixel = 91;
			1810: Pixel = 81;
			1811: Pixel = 97;
			1812: Pixel = 97;
			1813: Pixel = 97;
			1814: Pixel = 98;
			1815: Pixel = 101;
			1816: Pixel = 85;
			1817: Pixel = 160;
			1818: Pixel = 190;
			1819: Pixel = 154;
			1820: Pixel = 142;
			1821: Pixel = 116;
			1822: Pixel = 107;
			1823: Pixel = 135;
			1824: Pixel = 136;
			1825: Pixel = 122;
			1826: Pixel = 135;
			1827: Pixel = 146;
			1828: Pixel = 133;
			1829: Pixel = 141;
			1830: Pixel = 144;
			1831: Pixel = 154;
			1832: Pixel = 152;
			1833: Pixel = 153;
			1834: Pixel = 157;
			1835: Pixel = 143;
			1836: Pixel = 147;
			1837: Pixel = 161;
			1838: Pixel = 164;
			1839: Pixel = 165;
			1840: Pixel = 169;
			1841: Pixel = 168;
			1842: Pixel = 167;
			1843: Pixel = 159;
			1844: Pixel = 160;
			1845: Pixel = 170;
			1846: Pixel = 184;
			1847: Pixel = 193;
			1848: Pixel = 193;
			1849: Pixel = 191;
			1850: Pixel = 192;
			1851: Pixel = 195;
			1852: Pixel = 200;
			1853: Pixel = 201;
			1854: Pixel = 201;
			1855: Pixel = 212;
			1856: Pixel = 176;
			1857: Pixel = 151;
			1858: Pixel = 144;
			1859: Pixel = 179;
			1860: Pixel = 47;
			1861: Pixel = 48;
			1862: Pixel = 52;
			1863: Pixel = 51;
			1864: Pixel = 63;
			1865: Pixel = 142;
			1866: Pixel = 149;
			1867: Pixel = 157;
			1868: Pixel = 159;
			1869: Pixel = 156;
			1870: Pixel = 157;
			1871: Pixel = 157;
			1872: Pixel = 156;
			1873: Pixel = 156;
			1874: Pixel = 156;
			1875: Pixel = 98;
			1876: Pixel = 97;
			1877: Pixel = 98;
			1878: Pixel = 108;
			1879: Pixel = 140;
			1880: Pixel = 167;
			1881: Pixel = 173;
			1882: Pixel = 172;
			1883: Pixel = 149;
			1884: Pixel = 88;
			1885: Pixel = 78;
			1886: Pixel = 96;
			1887: Pixel = 97;
			1888: Pixel = 97;
			1889: Pixel = 98;
			1890: Pixel = 101;
			1891: Pixel = 82;
			1892: Pixel = 165;
			1893: Pixel = 201;
			1894: Pixel = 162;
			1895: Pixel = 155;
			1896: Pixel = 130;
			1897: Pixel = 118;
			1898: Pixel = 131;
			1899: Pixel = 120;
			1900: Pixel = 133;
			1901: Pixel = 141;
			1902: Pixel = 128;
			1903: Pixel = 133;
			1904: Pixel = 138;
			1905: Pixel = 147;
			1906: Pixel = 137;
			1907: Pixel = 125;
			1908: Pixel = 111;
			1909: Pixel = 106;
			1910: Pixel = 148;
			1911: Pixel = 133;
			1912: Pixel = 136;
			1913: Pixel = 141;
			1914: Pixel = 143;
			1915: Pixel = 140;
			1916: Pixel = 117;
			1917: Pixel = 115;
			1918: Pixel = 160;
			1919: Pixel = 170;
			1920: Pixel = 188;
			1921: Pixel = 197;
			1922: Pixel = 195;
			1923: Pixel = 190;
			1924: Pixel = 193;
			1925: Pixel = 199;
			1926: Pixel = 200;
			1927: Pixel = 202;
			1928: Pixel = 207;
			1929: Pixel = 217;
			1930: Pixel = 191;
			1931: Pixel = 124;
			1932: Pixel = 86;
			1933: Pixel = 175;
			1934: Pixel = 133;
			1935: Pixel = 28;
			1936: Pixel = 50;
			1937: Pixel = 51;
			1938: Pixel = 49;
			1939: Pixel = 100;
			1940: Pixel = 153;
			1941: Pixel = 151;
			1942: Pixel = 160;
			1943: Pixel = 157;
			1944: Pixel = 156;
			1945: Pixel = 156;
			1946: Pixel = 155;
			1947: Pixel = 155;
			1948: Pixel = 155;
			1949: Pixel = 153;
			1950: Pixel = 99;
			1951: Pixel = 99;
			1952: Pixel = 100;
			1953: Pixel = 111;
			1954: Pixel = 143;
			1955: Pixel = 169;
			1956: Pixel = 173;
			1957: Pixel = 173;
			1958: Pixel = 150;
			1959: Pixel = 89;
			1960: Pixel = 78;
			1961: Pixel = 95;
			1962: Pixel = 98;
			1963: Pixel = 99;
			1964: Pixel = 99;
			1965: Pixel = 102;
			1966: Pixel = 82;
			1967: Pixel = 153;
			1968: Pixel = 210;
			1969: Pixel = 170;
			1970: Pixel = 134;
			1971: Pixel = 127;
			1972: Pixel = 116;
			1973: Pixel = 114;
			1974: Pixel = 127;
			1975: Pixel = 138;
			1976: Pixel = 126;
			1977: Pixel = 130;
			1978: Pixel = 131;
			1979: Pixel = 139;
			1980: Pixel = 131;
			1981: Pixel = 130;
			1982: Pixel = 120;
			1983: Pixel = 105;
			1984: Pixel = 81;
			1985: Pixel = 123;
			1986: Pixel = 125;
			1987: Pixel = 81;
			1988: Pixel = 85;
			1989: Pixel = 77;
			1990: Pixel = 48;
			1991: Pixel = 39;
			1992: Pixel = 106;
			1993: Pixel = 174;
			1994: Pixel = 189;
			1995: Pixel = 197;
			1996: Pixel = 194;
			1997: Pixel = 194;
			1998: Pixel = 193;
			1999: Pixel = 196;
			2000: Pixel = 198;
			2001: Pixel = 204;
			2002: Pixel = 210;
			2003: Pixel = 183;
			2004: Pixel = 138;
			2005: Pixel = 96;
			2006: Pixel = 82;
			2007: Pixel = 152;
			2008: Pixel = 181;
			2009: Pixel = 48;
			2010: Pixel = 47;
			2011: Pixel = 49;
			2012: Pixel = 47;
			2013: Pixel = 53;
			2014: Pixel = 137;
			2015: Pixel = 149;
			2016: Pixel = 159;
			2017: Pixel = 160;
			2018: Pixel = 159;
			2019: Pixel = 157;
			2020: Pixel = 155;
			2021: Pixel = 154;
			2022: Pixel = 154;
			2023: Pixel = 153;
			2024: Pixel = 153;
			2025: Pixel = 103;
			2026: Pixel = 100;
			2027: Pixel = 99;
			2028: Pixel = 111;
			2029: Pixel = 142;
			2030: Pixel = 168;
			2031: Pixel = 171;
			2032: Pixel = 172;
			2033: Pixel = 150;
			2034: Pixel = 89;
			2035: Pixel = 79;
			2036: Pixel = 95;
			2037: Pixel = 97;
			2038: Pixel = 99;
			2039: Pixel = 99;
			2040: Pixel = 101;
			2041: Pixel = 85;
			2042: Pixel = 127;
			2043: Pixel = 214;
			2044: Pixel = 174;
			2045: Pixel = 127;
			2046: Pixel = 138;
			2047: Pixel = 110;
			2048: Pixel = 120;
			2049: Pixel = 138;
			2050: Pixel = 124;
			2051: Pixel = 128;
			2052: Pixel = 131;
			2053: Pixel = 136;
			2054: Pixel = 128;
			2055: Pixel = 128;
			2056: Pixel = 114;
			2057: Pixel = 100;
			2058: Pixel = 79;
			2059: Pixel = 61;
			2060: Pixel = 97;
			2061: Pixel = 84;
			2062: Pixel = 92;
			2063: Pixel = 81;
			2064: Pixel = 59;
			2065: Pixel = 41;
			2066: Pixel = 115;
			2067: Pixel = 166;
			2068: Pixel = 185;
			2069: Pixel = 194;
			2070: Pixel = 192;
			2071: Pixel = 189;
			2072: Pixel = 192;
			2073: Pixel = 191;
			2074: Pixel = 197;
			2075: Pixel = 207;
			2076: Pixel = 189;
			2077: Pixel = 146;
			2078: Pixel = 86;
			2079: Pixel = 89;
			2080: Pixel = 116;
			2081: Pixel = 173;
			2082: Pixel = 168;
			2083: Pixel = 47;
			2084: Pixel = 46;
			2085: Pixel = 49;
			2086: Pixel = 50;
			2087: Pixel = 49;
			2088: Pixel = 87;
			2089: Pixel = 151;
			2090: Pixel = 154;
			2091: Pixel = 164;
			2092: Pixel = 160;
			2093: Pixel = 160;
			2094: Pixel = 158;
			2095: Pixel = 156;
			2096: Pixel = 155;
			2097: Pixel = 154;
			2098: Pixel = 154;
			2099: Pixel = 152;
			2100: Pixel = 106;
			2101: Pixel = 103;
			2102: Pixel = 100;
			2103: Pixel = 108;
			2104: Pixel = 141;
			2105: Pixel = 167;
			2106: Pixel = 171;
			2107: Pixel = 171;
			2108: Pixel = 151;
			2109: Pixel = 91;
			2110: Pixel = 78;
			2111: Pixel = 94;
			2112: Pixel = 97;
			2113: Pixel = 99;
			2114: Pixel = 98;
			2115: Pixel = 99;
			2116: Pixel = 96;
			2117: Pixel = 99;
			2118: Pixel = 201;
			2119: Pixel = 188;
			2120: Pixel = 152;
			2121: Pixel = 132;
			2122: Pixel = 115;
			2123: Pixel = 137;
			2124: Pixel = 118;
			2125: Pixel = 124;
			2126: Pixel = 127;
			2127: Pixel = 125;
			2128: Pixel = 132;
			2129: Pixel = 126;
			2130: Pixel = 95;
			2131: Pixel = 73;
			2132: Pixel = 63;
			2133: Pixel = 44;
			2134: Pixel = 77;
			2135: Pixel = 90;
			2136: Pixel = 71;
			2137: Pixel = 91;
			2138: Pixel = 53;
			2139: Pixel = 76;
			2140: Pixel = 123;
			2141: Pixel = 170;
			2142: Pixel = 187;
			2143: Pixel = 181;
			2144: Pixel = 183;
			2145: Pixel = 183;
			2146: Pixel = 185;
			2147: Pixel = 189;
			2148: Pixel = 195;
			2149: Pixel = 189;
			2150: Pixel = 133;
			2151: Pixel = 101;
			2152: Pixel = 127;
			2153: Pixel = 147;
			2154: Pixel = 158;
			2155: Pixel = 189;
			2156: Pixel = 168;
			2157: Pixel = 46;
			2158: Pixel = 45;
			2159: Pixel = 56;
			2160: Pixel = 47;
			2161: Pixel = 50;
			2162: Pixel = 53;
			2163: Pixel = 128;
			2164: Pixel = 151;
			2165: Pixel = 162;
			2166: Pixel = 165;
			2167: Pixel = 163;
			2168: Pixel = 161;
			2169: Pixel = 158;
			2170: Pixel = 157;
			2171: Pixel = 155;
			2172: Pixel = 155;
			2173: Pixel = 154;
			2174: Pixel = 152;
			2175: Pixel = 107;
			2176: Pixel = 104;
			2177: Pixel = 99;
			2178: Pixel = 104;
			2179: Pixel = 139;
			2180: Pixel = 168;
			2181: Pixel = 171;
			2182: Pixel = 171;
			2183: Pixel = 152;
			2184: Pixel = 91;
			2185: Pixel = 77;
			2186: Pixel = 94;
			2187: Pixel = 96;
			2188: Pixel = 97;
			2189: Pixel = 97;
			2190: Pixel = 98;
			2191: Pixel = 105;
			2192: Pixel = 88;
			2193: Pixel = 168;
			2194: Pixel = 202;
			2195: Pixel = 169;
			2196: Pixel = 123;
			2197: Pixel = 129;
			2198: Pixel = 122;
			2199: Pixel = 123;
			2200: Pixel = 123;
			2201: Pixel = 124;
			2202: Pixel = 132;
			2203: Pixel = 97;
			2204: Pixel = 81;
			2205: Pixel = 73;
			2206: Pixel = 62;
			2207: Pixel = 65;
			2208: Pixel = 50;
			2209: Pixel = 76;
			2210: Pixel = 50;
			2211: Pixel = 83;
			2212: Pixel = 80;
			2213: Pixel = 74;
			2214: Pixel = 124;
			2215: Pixel = 170;
			2216: Pixel = 195;
			2217: Pixel = 184;
			2218: Pixel = 180;
			2219: Pixel = 178;
			2220: Pixel = 176;
			2221: Pixel = 184;
			2222: Pixel = 190;
			2223: Pixel = 186;
			2224: Pixel = 93;
			2225: Pixel = 77;
			2226: Pixel = 117;
			2227: Pixel = 128;
			2228: Pixel = 165;
			2229: Pixel = 190;
			2230: Pixel = 151;
			2231: Pixel = 49;
			2232: Pixel = 41;
			2233: Pixel = 56;
			2234: Pixel = 54;
			2235: Pixel = 47;
			2236: Pixel = 47;
			2237: Pixel = 76;
			2238: Pixel = 140;
			2239: Pixel = 153;
			2240: Pixel = 167;
			2241: Pixel = 164;
			2242: Pixel = 163;
			2243: Pixel = 162;
			2244: Pixel = 159;
			2245: Pixel = 158;
			2246: Pixel = 157;
			2247: Pixel = 156;
			2248: Pixel = 154;
			2249: Pixel = 152;
			2250: Pixel = 108;
			2251: Pixel = 105;
			2252: Pixel = 99;
			2253: Pixel = 98;
			2254: Pixel = 136;
			2255: Pixel = 168;
			2256: Pixel = 173;
			2257: Pixel = 173;
			2258: Pixel = 153;
			2259: Pixel = 90;
			2260: Pixel = 75;
			2261: Pixel = 92;
			2262: Pixel = 96;
			2263: Pixel = 96;
			2264: Pixel = 98;
			2265: Pixel = 100;
			2266: Pixel = 108;
			2267: Pixel = 102;
			2268: Pixel = 106;
			2269: Pixel = 200;
			2270: Pixel = 182;
			2271: Pixel = 131;
			2272: Pixel = 119;
			2273: Pixel = 122;
			2274: Pixel = 125;
			2275: Pixel = 122;
			2276: Pixel = 130;
			2277: Pixel = 108;
			2278: Pixel = 79;
			2279: Pixel = 84;
			2280: Pixel = 66;
			2281: Pixel = 51;
			2282: Pixel = 78;
			2283: Pixel = 53;
			2284: Pixel = 58;
			2285: Pixel = 62;
			2286: Pixel = 63;
			2287: Pixel = 82;
			2288: Pixel = 115;
			2289: Pixel = 147;
			2290: Pixel = 193;
			2291: Pixel = 186;
			2292: Pixel = 177;
			2293: Pixel = 178;
			2294: Pixel = 174;
			2295: Pixel = 178;
			2296: Pixel = 185;
			2297: Pixel = 189;
			2298: Pixel = 194;
			2299: Pixel = 122;
			2300: Pixel = 89;
			2301: Pixel = 106;
			2302: Pixel = 124;
			2303: Pixel = 163;
			2304: Pixel = 122;
			2305: Pixel = 37;
			2306: Pixel = 43;
			2307: Pixel = 56;
			2308: Pixel = 55;
			2309: Pixel = 49;
			2310: Pixel = 48;
			2311: Pixel = 52;
			2312: Pixel = 107;
			2313: Pixel = 133;
			2314: Pixel = 162;
			2315: Pixel = 166;
			2316: Pixel = 162;
			2317: Pixel = 163;
			2318: Pixel = 162;
			2319: Pixel = 161;
			2320: Pixel = 160;
			2321: Pixel = 159;
			2322: Pixel = 156;
			2323: Pixel = 155;
			2324: Pixel = 152;
			2325: Pixel = 106;
			2326: Pixel = 104;
			2327: Pixel = 98;
			2328: Pixel = 93;
			2329: Pixel = 133;
			2330: Pixel = 167;
			2331: Pixel = 173;
			2332: Pixel = 174;
			2333: Pixel = 154;
			2334: Pixel = 91;
			2335: Pixel = 74;
			2336: Pixel = 93;
			2337: Pixel = 98;
			2338: Pixel = 98;
			2339: Pixel = 97;
			2340: Pixel = 100;
			2341: Pixel = 109;
			2342: Pixel = 112;
			2343: Pixel = 94;
			2344: Pixel = 194;
			2345: Pixel = 194;
			2346: Pixel = 120;
			2347: Pixel = 116;
			2348: Pixel = 118;
			2349: Pixel = 128;
			2350: Pixel = 130;
			2351: Pixel = 102;
			2352: Pixel = 80;
			2353: Pixel = 52;
			2354: Pixel = 71;
			2355: Pixel = 74;
			2356: Pixel = 55;
			2357: Pixel = 84;
			2358: Pixel = 66;
			2359: Pixel = 46;
			2360: Pixel = 42;
			2361: Pixel = 63;
			2362: Pixel = 94;
			2363: Pixel = 135;
			2364: Pixel = 178;
			2365: Pixel = 182;
			2366: Pixel = 170;
			2367: Pixel = 172;
			2368: Pixel = 173;
			2369: Pixel = 170;
			2370: Pixel = 185;
			2371: Pixel = 197;
			2372: Pixel = 195;
			2373: Pixel = 203;
			2374: Pixel = 165;
			2375: Pixel = 74;
			2376: Pixel = 67;
			2377: Pixel = 119;
			2378: Pixel = 145;
			2379: Pixel = 52;
			2380: Pixel = 40;
			2381: Pixel = 54;
			2382: Pixel = 58;
			2383: Pixel = 57;
			2384: Pixel = 45;
			2385: Pixel = 45;
			2386: Pixel = 68;
			2387: Pixel = 127;
			2388: Pixel = 137;
			2389: Pixel = 165;
			2390: Pixel = 166;
			2391: Pixel = 164;
			2392: Pixel = 162;
			2393: Pixel = 162;
			2394: Pixel = 161;
			2395: Pixel = 160;
			2396: Pixel = 158;
			2397: Pixel = 157;
			2398: Pixel = 156;
			2399: Pixel = 152;
			2400: Pixel = 104;
			2401: Pixel = 104;
			2402: Pixel = 99;
			2403: Pixel = 94;
			2404: Pixel = 133;
			2405: Pixel = 166;
			2406: Pixel = 173;
			2407: Pixel = 173;
			2408: Pixel = 154;
			2409: Pixel = 93;
			2410: Pixel = 75;
			2411: Pixel = 94;
			2412: Pixel = 99;
			2413: Pixel = 101;
			2414: Pixel = 99;
			2415: Pixel = 102;
			2416: Pixel = 112;
			2417: Pixel = 115;
			2418: Pixel = 97;
			2419: Pixel = 190;
			2420: Pixel = 162;
			2421: Pixel = 100;
			2422: Pixel = 117;
			2423: Pixel = 121;
			2424: Pixel = 118;
			2425: Pixel = 109;
			2426: Pixel = 63;
			2427: Pixel = 60;
			2428: Pixel = 45;
			2429: Pixel = 53;
			2430: Pixel = 73;
			2431: Pixel = 64;
			2432: Pixel = 68;
			2433: Pixel = 90;
			2434: Pixel = 37;
			2435: Pixel = 52;
			2436: Pixel = 122;
			2437: Pixel = 148;
			2438: Pixel = 160;
			2439: Pixel = 185;
			2440: Pixel = 181;
			2441: Pixel = 163;
			2442: Pixel = 172;
			2443: Pixel = 165;
			2444: Pixel = 178;
			2445: Pixel = 196;
			2446: Pixel = 200;
			2447: Pixel = 200;
			2448: Pixel = 208;
			2449: Pixel = 185;
			2450: Pixel = 88;
			2451: Pixel = 41;
			2452: Pixel = 100;
			2453: Pixel = 146;
			2454: Pixel = 52;
			2455: Pixel = 48;
			2456: Pixel = 53;
			2457: Pixel = 60;
			2458: Pixel = 53;
			2459: Pixel = 47;
			2460: Pixel = 44;
			2461: Pixel = 97;
			2462: Pixel = 139;
			2463: Pixel = 147;
			2464: Pixel = 154;
			2465: Pixel = 159;
			2466: Pixel = 162;
			2467: Pixel = 161;
			2468: Pixel = 162;
			2469: Pixel = 163;
			2470: Pixel = 160;
			2471: Pixel = 158;
			2472: Pixel = 158;
			2473: Pixel = 156;
			2474: Pixel = 152;
			2475: Pixel = 104;
			2476: Pixel = 102;
			2477: Pixel = 98;
			2478: Pixel = 94;
			2479: Pixel = 132;
			2480: Pixel = 166;
			2481: Pixel = 173;
			2482: Pixel = 174;
			2483: Pixel = 154;
			2484: Pixel = 96;
			2485: Pixel = 78;
			2486: Pixel = 96;
			2487: Pixel = 102;
			2488: Pixel = 103;
			2489: Pixel = 99;
			2490: Pixel = 104;
			2491: Pixel = 122;
			2492: Pixel = 117;
			2493: Pixel = 106;
			2494: Pixel = 152;
			2495: Pixel = 156;
			2496: Pixel = 106;
			2497: Pixel = 121;
			2498: Pixel = 132;
			2499: Pixel = 93;
			2500: Pixel = 57;
			2501: Pixel = 57;
			2502: Pixel = 63;
			2503: Pixel = 52;
			2504: Pixel = 53;
			2505: Pixel = 51;
			2506: Pixel = 69;
			2507: Pixel = 85;
			2508: Pixel = 78;
			2509: Pixel = 42;
			2510: Pixel = 124;
			2511: Pixel = 168;
			2512: Pixel = 175;
			2513: Pixel = 153;
			2514: Pixel = 184;
			2515: Pixel = 174;
			2516: Pixel = 163;
			2517: Pixel = 158;
			2518: Pixel = 170;
			2519: Pixel = 189;
			2520: Pixel = 197;
			2521: Pixel = 201;
			2522: Pixel = 205;
			2523: Pixel = 212;
			2524: Pixel = 203;
			2525: Pixel = 115;
			2526: Pixel = 37;
			2527: Pixel = 69;
			2528: Pixel = 147;
			2529: Pixel = 60;
			2530: Pixel = 51;
			2531: Pixel = 58;
			2532: Pixel = 63;
			2533: Pixel = 50;
			2534: Pixel = 49;
			2535: Pixel = 51;
			2536: Pixel = 124;
			2537: Pixel = 146;
			2538: Pixel = 161;
			2539: Pixel = 152;
			2540: Pixel = 149;
			2541: Pixel = 149;
			2542: Pixel = 152;
			2543: Pixel = 154;
			2544: Pixel = 158;
			2545: Pixel = 160;
			2546: Pixel = 158;
			2547: Pixel = 156;
			2548: Pixel = 154;
			2549: Pixel = 151;
			2550: Pixel = 103;
			2551: Pixel = 101;
			2552: Pixel = 96;
			2553: Pixel = 92;
			2554: Pixel = 131;
			2555: Pixel = 167;
			2556: Pixel = 174;
			2557: Pixel = 174;
			2558: Pixel = 154;
			2559: Pixel = 94;
			2560: Pixel = 81;
			2561: Pixel = 97;
			2562: Pixel = 101;
			2563: Pixel = 103;
			2564: Pixel = 102;
			2565: Pixel = 106;
			2566: Pixel = 114;
			2567: Pixel = 117;
			2568: Pixel = 113;
			2569: Pixel = 124;
			2570: Pixel = 139;
			2571: Pixel = 119;
			2572: Pixel = 136;
			2573: Pixel = 105;
			2574: Pixel = 58;
			2575: Pixel = 64;
			2576: Pixel = 46;
			2577: Pixel = 64;
			2578: Pixel = 64;
			2579: Pixel = 48;
			2580: Pixel = 59;
			2581: Pixel = 59;
			2582: Pixel = 63;
			2583: Pixel = 63;
			2584: Pixel = 115;
			2585: Pixel = 152;
			2586: Pixel = 175;
			2587: Pixel = 182;
			2588: Pixel = 161;
			2589: Pixel = 185;
			2590: Pixel = 163;
			2591: Pixel = 158;
			2592: Pixel = 166;
			2593: Pixel = 175;
			2594: Pixel = 188;
			2595: Pixel = 197;
			2596: Pixel = 201;
			2597: Pixel = 205;
			2598: Pixel = 209;
			2599: Pixel = 211;
			2600: Pixel = 142;
			2601: Pixel = 54;
			2602: Pixel = 50;
			2603: Pixel = 141;
			2604: Pixel = 68;
			2605: Pixel = 50;
			2606: Pixel = 61;
			2607: Pixel = 59;
			2608: Pixel = 51;
			2609: Pixel = 45;
			2610: Pixel = 78;
			2611: Pixel = 141;
			2612: Pixel = 152;
			2613: Pixel = 165;
			2614: Pixel = 160;
			2615: Pixel = 159;
			2616: Pixel = 156;
			2617: Pixel = 151;
			2618: Pixel = 145;
			2619: Pixel = 146;
			2620: Pixel = 147;
			2621: Pixel = 149;
			2622: Pixel = 151;
			2623: Pixel = 153;
			2624: Pixel = 152;
			2625: Pixel = 101;
			2626: Pixel = 99;
			2627: Pixel = 97;
			2628: Pixel = 92;
			2629: Pixel = 132;
			2630: Pixel = 167;
			2631: Pixel = 175;
			2632: Pixel = 175;
			2633: Pixel = 154;
			2634: Pixel = 94;
			2635: Pixel = 78;
			2636: Pixel = 96;
			2637: Pixel = 102;
			2638: Pixel = 103;
			2639: Pixel = 102;
			2640: Pixel = 106;
			2641: Pixel = 116;
			2642: Pixel = 116;
			2643: Pixel = 128;
			2644: Pixel = 119;
			2645: Pixel = 110;
			2646: Pixel = 134;
			2647: Pixel = 121;
			2648: Pixel = 77;
			2649: Pixel = 55;
			2650: Pixel = 71;
			2651: Pixel = 48;
			2652: Pixel = 70;
			2653: Pixel = 55;
			2654: Pixel = 49;
			2655: Pixel = 59;
			2656: Pixel = 68;
			2657: Pixel = 51;
			2658: Pixel = 79;
			2659: Pixel = 148;
			2660: Pixel = 170;
			2661: Pixel = 162;
			2662: Pixel = 193;
			2663: Pixel = 168;
			2664: Pixel = 130;
			2665: Pixel = 144;
			2666: Pixel = 165;
			2667: Pixel = 182;
			2668: Pixel = 178;
			2669: Pixel = 181;
			2670: Pixel = 194;
			2671: Pixel = 195;
			2672: Pixel = 199;
			2673: Pixel = 209;
			2674: Pixel = 218;
			2675: Pixel = 153;
			2676: Pixel = 53;
			2677: Pixel = 39;
			2678: Pixel = 131;
			2679: Pixel = 86;
			2680: Pixel = 54;
			2681: Pixel = 64;
			2682: Pixel = 56;
			2683: Pixel = 51;
			2684: Pixel = 46;
			2685: Pixel = 110;
			2686: Pixel = 141;
			2687: Pixel = 158;
			2688: Pixel = 161;
			2689: Pixel = 159;
			2690: Pixel = 163;
			2691: Pixel = 165;
			2692: Pixel = 159;
			2693: Pixel = 153;
			2694: Pixel = 148;
			2695: Pixel = 144;
			2696: Pixel = 142;
			2697: Pixel = 142;
			2698: Pixel = 145;
			2699: Pixel = 147;
			2700: Pixel = 101;
			2701: Pixel = 101;
			2702: Pixel = 99;
			2703: Pixel = 92;
			2704: Pixel = 130;
			2705: Pixel = 167;
			2706: Pixel = 175;
			2707: Pixel = 176;
			2708: Pixel = 156;
			2709: Pixel = 95;
			2710: Pixel = 80;
			2711: Pixel = 96;
			2712: Pixel = 103;
			2713: Pixel = 101;
			2714: Pixel = 101;
			2715: Pixel = 106;
			2716: Pixel = 112;
			2717: Pixel = 120;
			2718: Pixel = 154;
			2719: Pixel = 68;
			2720: Pixel = 75;
			2721: Pixel = 142;
			2722: Pixel = 72;
			2723: Pixel = 72;
			2724: Pixel = 66;
			2725: Pixel = 80;
			2726: Pixel = 46;
			2727: Pixel = 64;
			2728: Pixel = 50;
			2729: Pixel = 44;
			2730: Pixel = 74;
			2731: Pixel = 60;
			2732: Pixel = 65;
			2733: Pixel = 140;
			2734: Pixel = 178;
			2735: Pixel = 174;
			2736: Pixel = 177;
			2737: Pixel = 182;
			2738: Pixel = 137;
			2739: Pixel = 132;
			2740: Pixel = 117;
			2741: Pixel = 94;
			2742: Pixel = 132;
			2743: Pixel = 174;
			2744: Pixel = 174;
			2745: Pixel = 189;
			2746: Pixel = 189;
			2747: Pixel = 195;
			2748: Pixel = 187;
			2749: Pixel = 150;
			2750: Pixel = 109;
			2751: Pixel = 59;
			2752: Pixel = 35;
			2753: Pixel = 119;
			2754: Pixel = 101;
			2755: Pixel = 54;
			2756: Pixel = 65;
			2757: Pixel = 51;
			2758: Pixel = 51;
			2759: Pixel = 60;
			2760: Pixel = 127;
			2761: Pixel = 144;
			2762: Pixel = 162;
			2763: Pixel = 157;
			2764: Pixel = 157;
			2765: Pixel = 156;
			2766: Pixel = 159;
			2767: Pixel = 158;
			2768: Pixel = 154;
			2769: Pixel = 154;
			2770: Pixel = 154;
			2771: Pixel = 151;
			2772: Pixel = 144;
			2773: Pixel = 140;
			2774: Pixel = 134;
			2775: Pixel = 101;
			2776: Pixel = 103;
			2777: Pixel = 98;
			2778: Pixel = 89;
			2779: Pixel = 129;
			2780: Pixel = 167;
			2781: Pixel = 175;
			2782: Pixel = 176;
			2783: Pixel = 157;
			2784: Pixel = 97;
			2785: Pixel = 78;
			2786: Pixel = 96;
			2787: Pixel = 102;
			2788: Pixel = 100;
			2789: Pixel = 99;
			2790: Pixel = 99;
			2791: Pixel = 120;
			2792: Pixel = 145;
			2793: Pixel = 153;
			2794: Pixel = 136;
			2795: Pixel = 98;
			2796: Pixel = 71;
			2797: Pixel = 78;
			2798: Pixel = 84;
			2799: Pixel = 74;
			2800: Pixel = 64;
			2801: Pixel = 61;
			2802: Pixel = 50;
			2803: Pixel = 75;
			2804: Pixel = 42;
			2805: Pixel = 50;
			2806: Pixel = 47;
			2807: Pixel = 120;
			2808: Pixel = 173;
			2809: Pixel = 189;
			2810: Pixel = 188;
			2811: Pixel = 154;
			2812: Pixel = 92;
			2813: Pixel = 90;
			2814: Pixel = 90;
			2815: Pixel = 81;
			2816: Pixel = 91;
			2817: Pixel = 107;
			2818: Pixel = 140;
			2819: Pixel = 163;
			2820: Pixel = 185;
			2821: Pixel = 199;
			2822: Pixel = 173;
			2823: Pixel = 97;
			2824: Pixel = 63;
			2825: Pixel = 81;
			2826: Pixel = 72;
			2827: Pixel = 36;
			2828: Pixel = 110;
			2829: Pixel = 112;
			2830: Pixel = 54;
			2831: Pixel = 61;
			2832: Pixel = 50;
			2833: Pixel = 47;
			2834: Pixel = 80;
			2835: Pixel = 137;
			2836: Pixel = 150;
			2837: Pixel = 160;
			2838: Pixel = 155;
			2839: Pixel = 156;
			2840: Pixel = 154;
			2841: Pixel = 156;
			2842: Pixel = 156;
			2843: Pixel = 153;
			2844: Pixel = 153;
			2845: Pixel = 155;
			2846: Pixel = 154;
			2847: Pixel = 149;
			2848: Pixel = 144;
			2849: Pixel = 136;
			2850: Pixel = 97;
			2851: Pixel = 95;
			2852: Pixel = 91;
			2853: Pixel = 80;
			2854: Pixel = 126;
			2855: Pixel = 168;
			2856: Pixel = 177;
			2857: Pixel = 176;
			2858: Pixel = 155;
			2859: Pixel = 95;
			2860: Pixel = 76;
			2861: Pixel = 94;
			2862: Pixel = 98;
			2863: Pixel = 100;
			2864: Pixel = 90;
			2865: Pixel = 119;
			2866: Pixel = 171;
			2867: Pixel = 140;
			2868: Pixel = 153;
			2869: Pixel = 96;
			2870: Pixel = 49;
			2871: Pixel = 71;
			2872: Pixel = 75;
			2873: Pixel = 87;
			2874: Pixel = 84;
			2875: Pixel = 44;
			2876: Pixel = 71;
			2877: Pixel = 49;
			2878: Pixel = 57;
			2879: Pixel = 74;
			2880: Pixel = 34;
			2881: Pixel = 82;
			2882: Pixel = 165;
			2883: Pixel = 178;
			2884: Pixel = 204;
			2885: Pixel = 155;
			2886: Pixel = 55;
			2887: Pixel = 51;
			2888: Pixel = 41;
			2889: Pixel = 68;
			2890: Pixel = 110;
			2891: Pixel = 60;
			2892: Pixel = 123;
			2893: Pixel = 133;
			2894: Pixel = 150;
			2895: Pixel = 196;
			2896: Pixel = 190;
			2897: Pixel = 67;
			2898: Pixel = 61;
			2899: Pixel = 91;
			2900: Pixel = 47;
			2901: Pixel = 53;
			2902: Pixel = 38;
			2903: Pixel = 104;
			2904: Pixel = 119;
			2905: Pixel = 60;
			2906: Pixel = 54;
			2907: Pixel = 50;
			2908: Pixel = 45;
			2909: Pixel = 103;
			2910: Pixel = 146;
			2911: Pixel = 157;
			2912: Pixel = 156;
			2913: Pixel = 153;
			2914: Pixel = 153;
			2915: Pixel = 154;
			2916: Pixel = 154;
			2917: Pixel = 154;
			2918: Pixel = 153;
			2919: Pixel = 151;
			2920: Pixel = 150;
			2921: Pixel = 148;
			2922: Pixel = 142;
			2923: Pixel = 137;
			2924: Pixel = 133;
			2925: Pixel = 98;
			2926: Pixel = 96;
			2927: Pixel = 89;
			2928: Pixel = 76;
			2929: Pixel = 124;
			2930: Pixel = 169;
			2931: Pixel = 178;
			2932: Pixel = 179;
			2933: Pixel = 156;
			2934: Pixel = 97;
			2935: Pixel = 82;
			2936: Pixel = 100;
			2937: Pixel = 102;
			2938: Pixel = 103;
			2939: Pixel = 77;
			2940: Pixel = 90;
			2941: Pixel = 172;
			2942: Pixel = 177;
			2943: Pixel = 81;
			2944: Pixel = 48;
			2945: Pixel = 72;
			2946: Pixel = 66;
			2947: Pixel = 62;
			2948: Pixel = 100;
			2949: Pixel = 82;
			2950: Pixel = 39;
			2951: Pixel = 55;
			2952: Pixel = 63;
			2953: Pixel = 42;
			2954: Pixel = 41;
			2955: Pixel = 53;
			2956: Pixel = 127;
			2957: Pixel = 169;
			2958: Pixel = 198;
			2959: Pixel = 172;
			2960: Pixel = 111;
			2961: Pixel = 82;
			2962: Pixel = 82;
			2963: Pixel = 86;
			2964: Pixel = 130;
			2965: Pixel = 219;
			2966: Pixel = 121;
			2967: Pixel = 107;
			2968: Pixel = 125;
			2969: Pixel = 149;
			2970: Pixel = 211;
			2971: Pixel = 141;
			2972: Pixel = 73;
			2973: Pixel = 107;
			2974: Pixel = 153;
			2975: Pixel = 53;
			2976: Pixel = 46;
			2977: Pixel = 44;
			2978: Pixel = 101;
			2979: Pixel = 125;
			2980: Pixel = 67;
			2981: Pixel = 51;
			2982: Pixel = 50;
			2983: Pixel = 53;
			2984: Pixel = 128;
			2985: Pixel = 149;
			2986: Pixel = 158;
			2987: Pixel = 154;
			2988: Pixel = 152;
			2989: Pixel = 152;
			2990: Pixel = 152;
			2991: Pixel = 152;
			2992: Pixel = 152;
			2993: Pixel = 150;
			2994: Pixel = 147;
			2995: Pixel = 145;
			2996: Pixel = 139;
			2997: Pixel = 130;
			2998: Pixel = 133;
			2999: Pixel = 150;
			3000: Pixel = 102;
			3001: Pixel = 99;
			3002: Pixel = 89;
			3003: Pixel = 75;
			3004: Pixel = 123;
			3005: Pixel = 168;
			3006: Pixel = 179;
			3007: Pixel = 182;
			3008: Pixel = 159;
			3009: Pixel = 101;
			3010: Pixel = 87;
			3011: Pixel = 104;
			3012: Pixel = 117;
			3013: Pixel = 85;
			3014: Pixel = 95;
			3015: Pixel = 139;
			3016: Pixel = 155;
			3017: Pixel = 85;
			3018: Pixel = 62;
			3019: Pixel = 95;
			3020: Pixel = 64;
			3021: Pixel = 63;
			3022: Pixel = 82;
			3023: Pixel = 108;
			3024: Pixel = 109;
			3025: Pixel = 54;
			3026: Pixel = 42;
			3027: Pixel = 49;
			3028: Pixel = 50;
			3029: Pixel = 33;
			3030: Pixel = 96;
			3031: Pixel = 161;
			3032: Pixel = 195;
			3033: Pixel = 169;
			3034: Pixel = 114;
			3035: Pixel = 137;
			3036: Pixel = 144;
			3037: Pixel = 121;
			3038: Pixel = 121;
			3039: Pixel = 147;
			3040: Pixel = 162;
			3041: Pixel = 155;
			3042: Pixel = 126;
			3043: Pixel = 124;
			3044: Pixel = 147;
			3045: Pixel = 212;
			3046: Pixel = 159;
			3047: Pixel = 130;
			3048: Pixel = 139;
			3049: Pixel = 102;
			3050: Pixel = 66;
			3051: Pixel = 53;
			3052: Pixel = 50;
			3053: Pixel = 95;
			3054: Pixel = 136;
			3055: Pixel = 66;
			3056: Pixel = 48;
			3057: Pixel = 48;
			3058: Pixel = 78;
			3059: Pixel = 138;
			3060: Pixel = 152;
			3061: Pixel = 156;
			3062: Pixel = 152;
			3063: Pixel = 150;
			3064: Pixel = 154;
			3065: Pixel = 152;
			3066: Pixel = 153;
			3067: Pixel = 150;
			3068: Pixel = 145;
			3069: Pixel = 142;
			3070: Pixel = 135;
			3071: Pixel = 136;
			3072: Pixel = 156;
			3073: Pixel = 178;
			3074: Pixel = 187;
			3075: Pixel = 100;
			3076: Pixel = 93;
			3077: Pixel = 83;
			3078: Pixel = 67;
			3079: Pixel = 119;
			3080: Pixel = 168;
			3081: Pixel = 179;
			3082: Pixel = 183;
			3083: Pixel = 162;
			3084: Pixel = 101;
			3085: Pixel = 85;
			3086: Pixel = 105;
			3087: Pixel = 105;
			3088: Pixel = 125;
			3089: Pixel = 143;
			3090: Pixel = 98;
			3091: Pixel = 68;
			3092: Pixel = 40;
			3093: Pixel = 80;
			3094: Pixel = 114;
			3095: Pixel = 68;
			3096: Pixel = 58;
			3097: Pixel = 86;
			3098: Pixel = 101;
			3099: Pixel = 112;
			3100: Pixel = 55;
			3101: Pixel = 44;
			3102: Pixel = 49;
			3103: Pixel = 41;
			3104: Pixel = 62;
			3105: Pixel = 137;
			3106: Pixel = 188;
			3107: Pixel = 173;
			3108: Pixel = 96;
			3109: Pixel = 130;
			3110: Pixel = 149;
			3111: Pixel = 154;
			3112: Pixel = 154;
			3113: Pixel = 144;
			3114: Pixel = 145;
			3115: Pixel = 156;
			3116: Pixel = 157;
			3117: Pixel = 134;
			3118: Pixel = 129;
			3119: Pixel = 139;
			3120: Pixel = 207;
			3121: Pixel = 190;
			3122: Pixel = 147;
			3123: Pixel = 127;
			3124: Pixel = 105;
			3125: Pixel = 97;
			3126: Pixel = 53;
			3127: Pixel = 49;
			3128: Pixel = 89;
			3129: Pixel = 146;
			3130: Pixel = 60;
			3131: Pixel = 49;
			3132: Pixel = 45;
			3133: Pixel = 99;
			3134: Pixel = 143;
			3135: Pixel = 155;
			3136: Pixel = 153;
			3137: Pixel = 151;
			3138: Pixel = 151;
			3139: Pixel = 150;
			3140: Pixel = 149;
			3141: Pixel = 149;
			3142: Pixel = 146;
			3143: Pixel = 142;
			3144: Pixel = 132;
			3145: Pixel = 144;
			3146: Pixel = 180;
			3147: Pixel = 193;
			3148: Pixel = 191;
			3149: Pixel = 188;
			3150: Pixel = 92;
			3151: Pixel = 86;
			3152: Pixel = 77;
			3153: Pixel = 61;
			3154: Pixel = 116;
			3155: Pixel = 167;
			3156: Pixel = 178;
			3157: Pixel = 182;
			3158: Pixel = 161;
			3159: Pixel = 101;
			3160: Pixel = 83;
			3161: Pixel = 104;
			3162: Pixel = 121;
			3163: Pixel = 135;
			3164: Pixel = 120;
			3165: Pixel = 93;
			3166: Pixel = 59;
			3167: Pixel = 78;
			3168: Pixel = 108;
			3169: Pixel = 93;
			3170: Pixel = 45;
			3171: Pixel = 54;
			3172: Pixel = 92;
			3173: Pixel = 106;
			3174: Pixel = 100;
			3175: Pixel = 77;
			3176: Pixel = 47;
			3177: Pixel = 47;
			3178: Pixel = 46;
			3179: Pixel = 106;
			3180: Pixel = 169;
			3181: Pixel = 189;
			3182: Pixel = 82;
			3183: Pixel = 109;
			3184: Pixel = 133;
			3185: Pixel = 149;
			3186: Pixel = 163;
			3187: Pixel = 172;
			3188: Pixel = 173;
			3189: Pixel = 174;
			3190: Pixel = 175;
			3191: Pixel = 158;
			3192: Pixel = 142;
			3193: Pixel = 131;
			3194: Pixel = 132;
			3195: Pixel = 201;
			3196: Pixel = 198;
			3197: Pixel = 160;
			3198: Pixel = 141;
			3199: Pixel = 131;
			3200: Pixel = 110;
			3201: Pixel = 57;
			3202: Pixel = 54;
			3203: Pixel = 79;
			3204: Pixel = 151;
			3205: Pixel = 55;
			3206: Pixel = 46;
			3207: Pixel = 49;
			3208: Pixel = 118;
			3209: Pixel = 147;
			3210: Pixel = 157;
			3211: Pixel = 152;
			3212: Pixel = 151;
			3213: Pixel = 151;
			3214: Pixel = 150;
			3215: Pixel = 147;
			3216: Pixel = 145;
			3217: Pixel = 142;
			3218: Pixel = 134;
			3219: Pixel = 144;
			3220: Pixel = 189;
			3221: Pixel = 199;
			3222: Pixel = 192;
			3223: Pixel = 188;
			3224: Pixel = 191;
			3225: Pixel = 83;
			3226: Pixel = 78;
			3227: Pixel = 73;
			3228: Pixel = 60;
			3229: Pixel = 116;
			3230: Pixel = 168;
			3231: Pixel = 177;
			3232: Pixel = 180;
			3233: Pixel = 160;
			3234: Pixel = 100;
			3235: Pixel = 81;
			3236: Pixel = 106;
			3237: Pixel = 121;
			3238: Pixel = 114;
			3239: Pixel = 89;
			3240: Pixel = 71;
			3241: Pixel = 73;
			3242: Pixel = 85;
			3243: Pixel = 111;
			3244: Pixel = 68;
			3245: Pixel = 44;
			3246: Pixel = 47;
			3247: Pixel = 62;
			3248: Pixel = 62;
			3249: Pixel = 63;
			3250: Pixel = 125;
			3251: Pixel = 48;
			3252: Pixel = 34;
			3253: Pixel = 70;
			3254: Pixel = 141;
			3255: Pixel = 200;
			3256: Pixel = 91;
			3257: Pixel = 66;
			3258: Pixel = 125;
			3259: Pixel = 129;
			3260: Pixel = 144;
			3261: Pixel = 158;
			3262: Pixel = 173;
			3263: Pixel = 179;
			3264: Pixel = 176;
			3265: Pixel = 171;
			3266: Pixel = 156;
			3267: Pixel = 146;
			3268: Pixel = 134;
			3269: Pixel = 130;
			3270: Pixel = 195;
			3271: Pixel = 201;
			3272: Pixel = 159;
			3273: Pixel = 144;
			3274: Pixel = 132;
			3275: Pixel = 109;
			3276: Pixel = 53;
			3277: Pixel = 58;
			3278: Pixel = 68;
			3279: Pixel = 153;
			3280: Pixel = 59;
			3281: Pixel = 44;
			3282: Pixel = 63;
			3283: Pixel = 136;
			3284: Pixel = 154;
			3285: Pixel = 156;
			3286: Pixel = 153;
			3287: Pixel = 150;
			3288: Pixel = 149;
			3289: Pixel = 148;
			3290: Pixel = 146;
			3291: Pixel = 144;
			3292: Pixel = 137;
			3293: Pixel = 134;
			3294: Pixel = 182;
			3295: Pixel = 197;
			3296: Pixel = 193;
			3297: Pixel = 193;
			3298: Pixel = 195;
			3299: Pixel = 201;
			3300: Pixel = 76;
			3301: Pixel = 75;
			3302: Pixel = 69;
			3303: Pixel = 55;
			3304: Pixel = 114;
			3305: Pixel = 166;
			3306: Pixel = 174;
			3307: Pixel = 175;
			3308: Pixel = 160;
			3309: Pixel = 99;
			3310: Pixel = 88;
			3311: Pixel = 105;
			3312: Pixel = 121;
			3313: Pixel = 101;
			3314: Pixel = 100;
			3315: Pixel = 97;
			3316: Pixel = 73;
			3317: Pixel = 75;
			3318: Pixel = 110;
			3319: Pixel = 62;
			3320: Pixel = 54;
			3321: Pixel = 44;
			3322: Pixel = 54;
			3323: Pixel = 52;
			3324: Pixel = 74;
			3325: Pixel = 130;
			3326: Pixel = 92;
			3327: Pixel = 31;
			3328: Pixel = 100;
			3329: Pixel = 188;
			3330: Pixel = 149;
			3331: Pixel = 34;
			3332: Pixel = 82;
			3333: Pixel = 120;
			3334: Pixel = 131;
			3335: Pixel = 141;
			3336: Pixel = 152;
			3337: Pixel = 164;
			3338: Pixel = 175;
			3339: Pixel = 173;
			3340: Pixel = 166;
			3341: Pixel = 148;
			3342: Pixel = 137;
			3343: Pixel = 129;
			3344: Pixel = 127;
			3345: Pixel = 184;
			3346: Pixel = 204;
			3347: Pixel = 156;
			3348: Pixel = 145;
			3349: Pixel = 135;
			3350: Pixel = 98;
			3351: Pixel = 47;
			3352: Pixel = 62;
			3353: Pixel = 58;
			3354: Pixel = 153;
			3355: Pixel = 76;
			3356: Pixel = 40;
			3357: Pixel = 87;
			3358: Pixel = 146;
			3359: Pixel = 160;
			3360: Pixel = 155;
			3361: Pixel = 153;
			3362: Pixel = 150;
			3363: Pixel = 147;
			3364: Pixel = 145;
			3365: Pixel = 143;
			3366: Pixel = 142;
			3367: Pixel = 130;
			3368: Pixel = 162;
			3369: Pixel = 197;
			3370: Pixel = 191;
			3371: Pixel = 193;
			3372: Pixel = 201;
			3373: Pixel = 206;
			3374: Pixel = 203;
			3375: Pixel = 78;
			3376: Pixel = 76;
			3377: Pixel = 66;
			3378: Pixel = 49;
			3379: Pixel = 112;
			3380: Pixel = 166;
			3381: Pixel = 173;
			3382: Pixel = 176;
			3383: Pixel = 160;
			3384: Pixel = 96;
			3385: Pixel = 81;
			3386: Pixel = 123;
			3387: Pixel = 130;
			3388: Pixel = 82;
			3389: Pixel = 99;
			3390: Pixel = 83;
			3391: Pixel = 79;
			3392: Pixel = 100;
			3393: Pixel = 121;
			3394: Pixel = 71;
			3395: Pixel = 48;
			3396: Pixel = 39;
			3397: Pixel = 68;
			3398: Pixel = 86;
			3399: Pixel = 114;
			3400: Pixel = 122;
			3401: Pixel = 55;
			3402: Pixel = 52;
			3403: Pixel = 141;
			3404: Pixel = 181;
			3405: Pixel = 46;
			3406: Pixel = 52;
			3407: Pixel = 81;
			3408: Pixel = 115;
			3409: Pixel = 129;
			3410: Pixel = 138;
			3411: Pixel = 150;
			3412: Pixel = 156;
			3413: Pixel = 162;
			3414: Pixel = 166;
			3415: Pixel = 162;
			3416: Pixel = 143;
			3417: Pixel = 129;
			3418: Pixel = 126;
			3419: Pixel = 122;
			3420: Pixel = 172;
			3421: Pixel = 212;
			3422: Pixel = 155;
			3423: Pixel = 143;
			3424: Pixel = 133;
			3425: Pixel = 79;
			3426: Pixel = 46;
			3427: Pixel = 70;
			3428: Pixel = 49;
			3429: Pixel = 147;
			3430: Pixel = 90;
			3431: Pixel = 35;
			3432: Pixel = 111;
			3433: Pixel = 151;
			3434: Pixel = 158;
			3435: Pixel = 153;
			3436: Pixel = 152;
			3437: Pixel = 151;
			3438: Pixel = 148;
			3439: Pixel = 146;
			3440: Pixel = 143;
			3441: Pixel = 135;
			3442: Pixel = 140;
			3443: Pixel = 190;
			3444: Pixel = 194;
			3445: Pixel = 193;
			3446: Pixel = 203;
			3447: Pixel = 208;
			3448: Pixel = 207;
			3449: Pixel = 204;
			3450: Pixel = 82;
			3451: Pixel = 77;
			3452: Pixel = 65;
			3453: Pixel = 44;
			3454: Pixel = 109;
			3455: Pixel = 166;
			3456: Pixel = 174;
			3457: Pixel = 178;
			3458: Pixel = 161;
			3459: Pixel = 100;
			3460: Pixel = 91;
			3461: Pixel = 113;
			3462: Pixel = 112;
			3463: Pixel = 79;
			3464: Pixel = 98;
			3465: Pixel = 77;
			3466: Pixel = 84;
			3467: Pixel = 81;
			3468: Pixel = 116;
			3469: Pixel = 74;
			3470: Pixel = 52;
			3471: Pixel = 44;
			3472: Pixel = 64;
			3473: Pixel = 95;
			3474: Pixel = 99;
			3475: Pixel = 44;
			3476: Pixel = 46;
			3477: Pixel = 129;
			3478: Pixel = 163;
			3479: Pixel = 103;
			3480: Pixel = 24;
			3481: Pixel = 69;
			3482: Pixel = 83;
			3483: Pixel = 114;
			3484: Pixel = 128;
			3485: Pixel = 135;
			3486: Pixel = 145;
			3487: Pixel = 150;
			3488: Pixel = 155;
			3489: Pixel = 160;
			3490: Pixel = 157;
			3491: Pixel = 132;
			3492: Pixel = 125;
			3493: Pixel = 135;
			3494: Pixel = 125;
			3495: Pixel = 161;
			3496: Pixel = 211;
			3497: Pixel = 151;
			3498: Pixel = 141;
			3499: Pixel = 123;
			3500: Pixel = 54;
			3501: Pixel = 49;
			3502: Pixel = 70;
			3503: Pixel = 41;
			3504: Pixel = 138;
			3505: Pixel = 109;
			3506: Pixel = 41;
			3507: Pixel = 135;
			3508: Pixel = 153;
			3509: Pixel = 156;
			3510: Pixel = 151;
			3511: Pixel = 150;
			3512: Pixel = 149;
			3513: Pixel = 148;
			3514: Pixel = 147;
			3515: Pixel = 143;
			3516: Pixel = 131;
			3517: Pixel = 165;
			3518: Pixel = 199;
			3519: Pixel = 192;
			3520: Pixel = 201;
			3521: Pixel = 208;
			3522: Pixel = 204;
			3523: Pixel = 206;
			3524: Pixel = 207;
			3525: Pixel = 81;
			3526: Pixel = 78;
			3527: Pixel = 68;
			3528: Pixel = 60;
			3529: Pixel = 121;
			3530: Pixel = 165;
			3531: Pixel = 172;
			3532: Pixel = 178;
			3533: Pixel = 162;
			3534: Pixel = 105;
			3535: Pixel = 85;
			3536: Pixel = 103;
			3537: Pixel = 104;
			3538: Pixel = 80;
			3539: Pixel = 96;
			3540: Pixel = 71;
			3541: Pixel = 93;
			3542: Pixel = 73;
			3543: Pixel = 119;
			3544: Pixel = 104;
			3545: Pixel = 51;
			3546: Pixel = 66;
			3547: Pixel = 40;
			3548: Pixel = 75;
			3549: Pixel = 69;
			3550: Pixel = 29;
			3551: Pixel = 93;
			3552: Pixel = 195;
			3553: Pixel = 137;
			3554: Pixel = 39;
			3555: Pixel = 41;
			3556: Pixel = 71;
			3557: Pixel = 93;
			3558: Pixel = 114;
			3559: Pixel = 126;
			3560: Pixel = 134;
			3561: Pixel = 143;
			3562: Pixel = 149;
			3563: Pixel = 152;
			3564: Pixel = 157;
			3565: Pixel = 157;
			3566: Pixel = 139;
			3567: Pixel = 123;
			3568: Pixel = 104;
			3569: Pixel = 105;
			3570: Pixel = 139;
			3571: Pixel = 182;
			3572: Pixel = 146;
			3573: Pixel = 141;
			3574: Pixel = 96;
			3575: Pixel = 40;
			3576: Pixel = 56;
			3577: Pixel = 69;
			3578: Pixel = 38;
			3579: Pixel = 122;
			3580: Pixel = 119;
			3581: Pixel = 65;
			3582: Pixel = 149;
			3583: Pixel = 155;
			3584: Pixel = 154;
			3585: Pixel = 150;
			3586: Pixel = 150;
			3587: Pixel = 148;
			3588: Pixel = 146;
			3589: Pixel = 145;
			3590: Pixel = 140;
			3591: Pixel = 135;
			3592: Pixel = 183;
			3593: Pixel = 197;
			3594: Pixel = 198;
			3595: Pixel = 206;
			3596: Pixel = 206;
			3597: Pixel = 208;
			3598: Pixel = 209;
			3599: Pixel = 207;
			3600: Pixel = 77;
			3601: Pixel = 78;
			3602: Pixel = 69;
			3603: Pixel = 79;
			3604: Pixel = 136;
			3605: Pixel = 165;
			3606: Pixel = 170;
			3607: Pixel = 178;
			3608: Pixel = 165;
			3609: Pixel = 103;
			3610: Pixel = 77;
			3611: Pixel = 103;
			3612: Pixel = 112;
			3613: Pixel = 66;
			3614: Pixel = 75;
			3615: Pixel = 82;
			3616: Pixel = 71;
			3617: Pixel = 90;
			3618: Pixel = 108;
			3619: Pixel = 127;
			3620: Pixel = 57;
			3621: Pixel = 97;
			3622: Pixel = 69;
			3623: Pixel = 59;
			3624: Pixel = 88;
			3625: Pixel = 131;
			3626: Pixel = 119;
			3627: Pixel = 151;
			3628: Pixel = 53;
			3629: Pixel = 52;
			3630: Pixel = 47;
			3631: Pixel = 76;
			3632: Pixel = 101;
			3633: Pixel = 117;
			3634: Pixel = 126;
			3635: Pixel = 132;
			3636: Pixel = 141;
			3637: Pixel = 145;
			3638: Pixel = 150;
			3639: Pixel = 155;
			3640: Pixel = 158;
			3641: Pixel = 153;
			3642: Pixel = 138;
			3643: Pixel = 139;
			3644: Pixel = 147;
			3645: Pixel = 178;
			3646: Pixel = 173;
			3647: Pixel = 145;
			3648: Pixel = 133;
			3649: Pixel = 63;
			3650: Pixel = 43;
			3651: Pixel = 64;
			3652: Pixel = 77;
			3653: Pixel = 43;
			3654: Pixel = 103;
			3655: Pixel = 125;
			3656: Pixel = 96;
			3657: Pixel = 153;
			3658: Pixel = 155;
			3659: Pixel = 153;
			3660: Pixel = 150;
			3661: Pixel = 148;
			3662: Pixel = 148;
			3663: Pixel = 146;
			3664: Pixel = 145;
			3665: Pixel = 136;
			3666: Pixel = 144;
			3667: Pixel = 192;
			3668: Pixel = 197;
			3669: Pixel = 206;
			3670: Pixel = 207;
			3671: Pixel = 206;
			3672: Pixel = 209;
			3673: Pixel = 209;
			3674: Pixel = 209;
			3675: Pixel = 74;
			3676: Pixel = 74;
			3677: Pixel = 65;
			3678: Pixel = 80;
			3679: Pixel = 139;
			3680: Pixel = 165;
			3681: Pixel = 170;
			3682: Pixel = 178;
			3683: Pixel = 165;
			3684: Pixel = 105;
			3685: Pixel = 74;
			3686: Pixel = 113;
			3687: Pixel = 116;
			3688: Pixel = 73;
			3689: Pixel = 95;
			3690: Pixel = 61;
			3691: Pixel = 60;
			3692: Pixel = 77;
			3693: Pixel = 88;
			3694: Pixel = 112;
			3695: Pixel = 114;
			3696: Pixel = 80;
			3697: Pixel = 53;
			3698: Pixel = 77;
			3699: Pixel = 171;
			3700: Pixel = 143;
			3701: Pixel = 116;
			3702: Pixel = 83;
			3703: Pixel = 41;
			3704: Pixel = 59;
			3705: Pixel = 52;
			3706: Pixel = 71;
			3707: Pixel = 104;
			3708: Pixel = 117;
			3709: Pixel = 127;
			3710: Pixel = 133;
			3711: Pixel = 140;
			3712: Pixel = 140;
			3713: Pixel = 146;
			3714: Pixel = 152;
			3715: Pixel = 153;
			3716: Pixel = 151;
			3717: Pixel = 148;
			3718: Pixel = 171;
			3719: Pixel = 198;
			3720: Pixel = 202;
			3721: Pixel = 173;
			3722: Pixel = 145;
			3723: Pixel = 107;
			3724: Pixel = 43;
			3725: Pixel = 49;
			3726: Pixel = 70;
			3727: Pixel = 75;
			3728: Pixel = 46;
			3729: Pixel = 85;
			3730: Pixel = 131;
			3731: Pixel = 121;
			3732: Pixel = 152;
			3733: Pixel = 155;
			3734: Pixel = 152;
			3735: Pixel = 149;
			3736: Pixel = 148;
			3737: Pixel = 145;
			3738: Pixel = 145;
			3739: Pixel = 145;
			3740: Pixel = 133;
			3741: Pixel = 153;
			3742: Pixel = 196;
			3743: Pixel = 201;
			3744: Pixel = 208;
			3745: Pixel = 206;
			3746: Pixel = 206;
			3747: Pixel = 209;
			3748: Pixel = 210;
			3749: Pixel = 211;
			3750: Pixel = 65;
			3751: Pixel = 67;
			3752: Pixel = 64;
			3753: Pixel = 77;
			3754: Pixel = 136;
			3755: Pixel = 166;
			3756: Pixel = 172;
			3757: Pixel = 179;
			3758: Pixel = 168;
			3759: Pixel = 99;
			3760: Pixel = 82;
			3761: Pixel = 118;
			3762: Pixel = 98;
			3763: Pixel = 78;
			3764: Pixel = 77;
			3765: Pixel = 57;
			3766: Pixel = 73;
			3767: Pixel = 82;
			3768: Pixel = 75;
			3769: Pixel = 79;
			3770: Pixel = 125;
			3771: Pixel = 74;
			3772: Pixel = 96;
			3773: Pixel = 165;
			3774: Pixel = 162;
			3775: Pixel = 111;
			3776: Pixel = 93;
			3777: Pixel = 47;
			3778: Pixel = 56;
			3779: Pixel = 55;
			3780: Pixel = 59;
			3781: Pixel = 63;
			3782: Pixel = 96;
			3783: Pixel = 110;
			3784: Pixel = 129;
			3785: Pixel = 131;
			3786: Pixel = 138;
			3787: Pixel = 139;
			3788: Pixel = 137;
			3789: Pixel = 134;
			3790: Pixel = 141;
			3791: Pixel = 142;
			3792: Pixel = 142;
			3793: Pixel = 152;
			3794: Pixel = 172;
			3795: Pixel = 170;
			3796: Pixel = 146;
			3797: Pixel = 138;
			3798: Pixel = 69;
			3799: Pixel = 45;
			3800: Pixel = 53;
			3801: Pixel = 71;
			3802: Pixel = 76;
			3803: Pixel = 48;
			3804: Pixel = 72;
			3805: Pixel = 135;
			3806: Pixel = 132;
			3807: Pixel = 152;
			3808: Pixel = 155;
			3809: Pixel = 150;
			3810: Pixel = 147;
			3811: Pixel = 148;
			3812: Pixel = 146;
			3813: Pixel = 144;
			3814: Pixel = 143;
			3815: Pixel = 130;
			3816: Pixel = 156;
			3817: Pixel = 201;
			3818: Pixel = 208;
			3819: Pixel = 208;
			3820: Pixel = 208;
			3821: Pixel = 208;
			3822: Pixel = 211;
			3823: Pixel = 212;
			3824: Pixel = 211;
			3825: Pixel = 56;
			3826: Pixel = 63;
			3827: Pixel = 63;
			3828: Pixel = 82;
			3829: Pixel = 139;
			3830: Pixel = 169;
			3831: Pixel = 176;
			3832: Pixel = 180;
			3833: Pixel = 163;
			3834: Pixel = 109;
			3835: Pixel = 101;
			3836: Pixel = 110;
			3837: Pixel = 110;
			3838: Pixel = 54;
			3839: Pixel = 61;
			3840: Pixel = 61;
			3841: Pixel = 74;
			3842: Pixel = 114;
			3843: Pixel = 91;
			3844: Pixel = 91;
			3845: Pixel = 86;
			3846: Pixel = 98;
			3847: Pixel = 150;
			3848: Pixel = 202;
			3849: Pixel = 116;
			3850: Pixel = 123;
			3851: Pixel = 48;
			3852: Pixel = 51;
			3853: Pixel = 52;
			3854: Pixel = 55;
			3855: Pixel = 62;
			3856: Pixel = 61;
			3857: Pixel = 84;
			3858: Pixel = 101;
			3859: Pixel = 127;
			3860: Pixel = 127;
			3861: Pixel = 133;
			3862: Pixel = 144;
			3863: Pixel = 138;
			3864: Pixel = 107;
			3865: Pixel = 108;
			3866: Pixel = 118;
			3867: Pixel = 117;
			3868: Pixel = 118;
			3869: Pixel = 137;
			3870: Pixel = 116;
			3871: Pixel = 129;
			3872: Pixel = 114;
			3873: Pixel = 43;
			3874: Pixel = 49;
			3875: Pixel = 55;
			3876: Pixel = 70;
			3877: Pixel = 74;
			3878: Pixel = 56;
			3879: Pixel = 62;
			3880: Pixel = 140;
			3881: Pixel = 144;
			3882: Pixel = 153;
			3883: Pixel = 154;
			3884: Pixel = 151;
			3885: Pixel = 149;
			3886: Pixel = 147;
			3887: Pixel = 146;
			3888: Pixel = 144;
			3889: Pixel = 144;
			3890: Pixel = 128;
			3891: Pixel = 162;
			3892: Pixel = 208;
			3893: Pixel = 211;
			3894: Pixel = 209;
			3895: Pixel = 208;
			3896: Pixel = 210;
			3897: Pixel = 212;
			3898: Pixel = 213;
			3899: Pixel = 213;
			3900: Pixel = 55;
			3901: Pixel = 59;
			3902: Pixel = 60;
			3903: Pixel = 87;
			3904: Pixel = 137;
			3905: Pixel = 168;
			3906: Pixel = 177;
			3907: Pixel = 181;
			3908: Pixel = 166;
			3909: Pixel = 122;
			3910: Pixel = 82;
			3911: Pixel = 123;
			3912: Pixel = 94;
			3913: Pixel = 78;
			3914: Pixel = 50;
			3915: Pixel = 68;
			3916: Pixel = 94;
			3917: Pixel = 110;
			3918: Pixel = 84;
			3919: Pixel = 98;
			3920: Pixel = 88;
			3921: Pixel = 133;
			3922: Pixel = 147;
			3923: Pixel = 146;
			3924: Pixel = 142;
			3925: Pixel = 76;
			3926: Pixel = 47;
			3927: Pixel = 49;
			3928: Pixel = 51;
			3929: Pixel = 55;
			3930: Pixel = 62;
			3931: Pixel = 61;
			3932: Pixel = 75;
			3933: Pixel = 90;
			3934: Pixel = 116;
			3935: Pixel = 121;
			3936: Pixel = 127;
			3937: Pixel = 137;
			3938: Pixel = 146;
			3939: Pixel = 137;
			3940: Pixel = 124;
			3941: Pixel = 124;
			3942: Pixel = 141;
			3943: Pixel = 162;
			3944: Pixel = 164;
			3945: Pixel = 148;
			3946: Pixel = 146;
			3947: Pixel = 62;
			3948: Pixel = 44;
			3949: Pixel = 49;
			3950: Pixel = 52;
			3951: Pixel = 71;
			3952: Pixel = 76;
			3953: Pixel = 64;
			3954: Pixel = 61;
			3955: Pixel = 146;
			3956: Pixel = 151;
			3957: Pixel = 153;
			3958: Pixel = 154;
			3959: Pixel = 153;
			3960: Pixel = 151;
			3961: Pixel = 148;
			3962: Pixel = 146;
			3963: Pixel = 145;
			3964: Pixel = 143;
			3965: Pixel = 126;
			3966: Pixel = 171;
			3967: Pixel = 216;
			3968: Pixel = 210;
			3969: Pixel = 210;
			3970: Pixel = 212;
			3971: Pixel = 213;
			3972: Pixel = 211;
			3973: Pixel = 208;
			3974: Pixel = 207;
			3975: Pixel = 52;
			3976: Pixel = 52;
			3977: Pixel = 57;
			3978: Pixel = 89;
			3979: Pixel = 129;
			3980: Pixel = 165;
			3981: Pixel = 178;
			3982: Pixel = 180;
			3983: Pixel = 168;
			3984: Pixel = 94;
			3985: Pixel = 88;
			3986: Pixel = 118;
			3987: Pixel = 72;
			3988: Pixel = 85;
			3989: Pixel = 54;
			3990: Pixel = 64;
			3991: Pixel = 108;
			3992: Pixel = 123;
			3993: Pixel = 98;
			3994: Pixel = 94;
			3995: Pixel = 121;
			3996: Pixel = 117;
			3997: Pixel = 150;
			3998: Pixel = 177;
			3999: Pixel = 94;
			4000: Pixel = 42;
			4001: Pixel = 58;
			4002: Pixel = 52;
			4003: Pixel = 53;
			4004: Pixel = 58;
			4005: Pixel = 62;
			4006: Pixel = 60;
			4007: Pixel = 70;
			4008: Pixel = 74;
			4009: Pixel = 102;
			4010: Pixel = 112;
			4011: Pixel = 123;
			4012: Pixel = 132;
			4013: Pixel = 139;
			4014: Pixel = 139;
			4015: Pixel = 131;
			4016: Pixel = 128;
			4017: Pixel = 126;
			4018: Pixel = 128;
			4019: Pixel = 134;
			4020: Pixel = 149;
			4021: Pixel = 99;
			4022: Pixel = 40;
			4023: Pixel = 49;
			4024: Pixel = 56;
			4025: Pixel = 51;
			4026: Pixel = 74;
			4027: Pixel = 78;
			4028: Pixel = 67;
			4029: Pixel = 62;
			4030: Pixel = 147;
			4031: Pixel = 153;
			4032: Pixel = 153;
			4033: Pixel = 154;
			4034: Pixel = 154;
			4035: Pixel = 153;
			4036: Pixel = 151;
			4037: Pixel = 147;
			4038: Pixel = 144;
			4039: Pixel = 140;
			4040: Pixel = 121;
			4041: Pixel = 175;
			4042: Pixel = 220;
			4043: Pixel = 212;
			4044: Pixel = 214;
			4045: Pixel = 215;
			4046: Pixel = 210;
			4047: Pixel = 206;
			4048: Pixel = 206;
			4049: Pixel = 206;
			4050: Pixel = 50;
			4051: Pixel = 46;
			4052: Pixel = 65;
			4053: Pixel = 104;
			4054: Pixel = 127;
			4055: Pixel = 162;
			4056: Pixel = 176;
			4057: Pixel = 178;
			4058: Pixel = 165;
			4059: Pixel = 99;
			4060: Pixel = 87;
			4061: Pixel = 104;
			4062: Pixel = 78;
			4063: Pixel = 66;
			4064: Pixel = 54;
			4065: Pixel = 57;
			4066: Pixel = 97;
			4067: Pixel = 117;
			4068: Pixel = 127;
			4069: Pixel = 100;
			4070: Pixel = 104;
			4071: Pixel = 97;
			4072: Pixel = 151;
			4073: Pixel = 133;
			4074: Pixel = 37;
			4075: Pixel = 53;
			4076: Pixel = 56;
			4077: Pixel = 51;
			4078: Pixel = 52;
			4079: Pixel = 51;
			4080: Pixel = 58;
			4081: Pixel = 55;
			4082: Pixel = 60;
			4083: Pixel = 63;
			4084: Pixel = 77;
			4085: Pixel = 102;
			4086: Pixel = 120;
			4087: Pixel = 132;
			4088: Pixel = 137;
			4089: Pixel = 140;
			4090: Pixel = 145;
			4091: Pixel = 150;
			4092: Pixel = 161;
			4093: Pixel = 161;
			4094: Pixel = 159;
			4095: Pixel = 134;
			4096: Pixel = 56;
			4097: Pixel = 45;
			4098: Pixel = 53;
			4099: Pixel = 59;
			4100: Pixel = 50;
			4101: Pixel = 81;
			4102: Pixel = 81;
			4103: Pixel = 71;
			4104: Pixel = 61;
			4105: Pixel = 148;
			4106: Pixel = 154;
			4107: Pixel = 155;
			4108: Pixel = 154;
			4109: Pixel = 152;
			4110: Pixel = 152;
			4111: Pixel = 151;
			4112: Pixel = 147;
			4113: Pixel = 142;
			4114: Pixel = 138;
			4115: Pixel = 118;
			4116: Pixel = 180;
			4117: Pixel = 223;
			4118: Pixel = 213;
			4119: Pixel = 213;
			4120: Pixel = 212;
			4121: Pixel = 210;
			4122: Pixel = 208;
			4123: Pixel = 209;
			4124: Pixel = 213;
			4125: Pixel = 49;
			4126: Pixel = 46;
			4127: Pixel = 65;
			4128: Pixel = 101;
			4129: Pixel = 131;
			4130: Pixel = 163;
			4131: Pixel = 176;
			4132: Pixel = 178;
			4133: Pixel = 167;
			4134: Pixel = 99;
			4135: Pixel = 74;
			4136: Pixel = 82;
			4137: Pixel = 71;
			4138: Pixel = 70;
			4139: Pixel = 58;
			4140: Pixel = 53;
			4141: Pixel = 94;
			4142: Pixel = 80;
			4143: Pixel = 98;
			4144: Pixel = 126;
			4145: Pixel = 120;
			4146: Pixel = 124;
			4147: Pixel = 96;
			4148: Pixel = 62;
			4149: Pixel = 51;
			4150: Pixel = 52;
			4151: Pixel = 59;
			4152: Pixel = 52;
			4153: Pixel = 53;
			4154: Pixel = 49;
			4155: Pixel = 52;
			4156: Pixel = 56;
			4157: Pixel = 57;
			4158: Pixel = 63;
			4159: Pixel = 57;
			4160: Pixel = 60;
			4161: Pixel = 94;
			4162: Pixel = 119;
			4163: Pixel = 131;
			4164: Pixel = 142;
			4165: Pixel = 152;
			4166: Pixel = 165;
			4167: Pixel = 168;
			4168: Pixel = 167;
			4169: Pixel = 162;
			4170: Pixel = 103;
			4171: Pixel = 49;
			4172: Pixel = 55;
			4173: Pixel = 58;
			4174: Pixel = 56;
			4175: Pixel = 52;
			4176: Pixel = 88;
			4177: Pixel = 82;
			4178: Pixel = 75;
			4179: Pixel = 65;
			4180: Pixel = 148;
			4181: Pixel = 155;
			4182: Pixel = 155;
			4183: Pixel = 153;
			4184: Pixel = 151;
			4185: Pixel = 150;
			4186: Pixel = 149;
			4187: Pixel = 144;
			4188: Pixel = 139;
			4189: Pixel = 135;
			4190: Pixel = 120;
			4191: Pixel = 193;
			4192: Pixel = 222;
			4193: Pixel = 210;
			4194: Pixel = 213;
			4195: Pixel = 214;
			4196: Pixel = 209;
			4197: Pixel = 212;
			4198: Pixel = 207;
			4199: Pixel = 180;
			4200: Pixel = 47;
			4201: Pixel = 44;
			4202: Pixel = 51;
			4203: Pixel = 92;
			4204: Pixel = 130;
			4205: Pixel = 164;
			4206: Pixel = 173;
			4207: Pixel = 178;
			4208: Pixel = 163;
			4209: Pixel = 97;
			4210: Pixel = 112;
			4211: Pixel = 85;
			4212: Pixel = 62;
			4213: Pixel = 69;
			4214: Pixel = 62;
			4215: Pixel = 40;
			4216: Pixel = 91;
			4217: Pixel = 116;
			4218: Pixel = 71;
			4219: Pixel = 107;
			4220: Pixel = 119;
			4221: Pixel = 141;
			4222: Pixel = 125;
			4223: Pixel = 80;
			4224: Pixel = 41;
			4225: Pixel = 55;
			4226: Pixel = 66;
			4227: Pixel = 53;
			4228: Pixel = 53;
			4229: Pixel = 51;
			4230: Pixel = 48;
			4231: Pixel = 55;
			4232: Pixel = 61;
			4233: Pixel = 59;
			4234: Pixel = 68;
			4235: Pixel = 60;
			4236: Pixel = 75;
			4237: Pixel = 96;
			4238: Pixel = 114;
			4239: Pixel = 128;
			4240: Pixel = 143;
			4241: Pixel = 156;
			4242: Pixel = 164;
			4243: Pixel = 158;
			4244: Pixel = 152;
			4245: Pixel = 95;
			4246: Pixel = 42;
			4247: Pixel = 50;
			4248: Pixel = 61;
			4249: Pixel = 57;
			4250: Pixel = 54;
			4251: Pixel = 90;
			4252: Pixel = 85;
			4253: Pixel = 80;
			4254: Pixel = 71;
			4255: Pixel = 150;
			4256: Pixel = 133;
			4257: Pixel = 125;
			4258: Pixel = 138;
			4259: Pixel = 143;
			4260: Pixel = 148;
			4261: Pixel = 149;
			4262: Pixel = 144;
			4263: Pixel = 139;
			4264: Pixel = 128;
			4265: Pixel = 127;
			4266: Pixel = 208;
			4267: Pixel = 217;
			4268: Pixel = 210;
			4269: Pixel = 211;
			4270: Pixel = 208;
			4271: Pixel = 201;
			4272: Pixel = 160;
			4273: Pixel = 88;
			4274: Pixel = 51;
			4275: Pixel = 57;
			4276: Pixel = 46;
			4277: Pixel = 46;
			4278: Pixel = 72;
			4279: Pixel = 118;
			4280: Pixel = 163;
			4281: Pixel = 172;
			4282: Pixel = 174;
			4283: Pixel = 159;
			4284: Pixel = 140;
			4285: Pixel = 102;
			4286: Pixel = 76;
			4287: Pixel = 56;
			4288: Pixel = 69;
			4289: Pixel = 63;
			4290: Pixel = 54;
			4291: Pixel = 73;
			4292: Pixel = 136;
			4293: Pixel = 78;
			4294: Pixel = 98;
			4295: Pixel = 113;
			4296: Pixel = 116;
			4297: Pixel = 102;
			4298: Pixel = 134;
			4299: Pixel = 81;
			4300: Pixel = 48;
			4301: Pixel = 69;
			4302: Pixel = 54;
			4303: Pixel = 54;
			4304: Pixel = 50;
			4305: Pixel = 49;
			4306: Pixel = 52;
			4307: Pixel = 59;
			4308: Pixel = 53;
			4309: Pixel = 63;
			4310: Pixel = 100;
			4311: Pixel = 125;
			4312: Pixel = 129;
			4313: Pixel = 134;
			4314: Pixel = 136;
			4315: Pixel = 146;
			4316: Pixel = 151;
			4317: Pixel = 149;
			4318: Pixel = 157;
			4319: Pixel = 179;
			4320: Pixel = 188;
			4321: Pixel = 150;
			4322: Pixel = 87;
			4323: Pixel = 47;
			4324: Pixel = 44;
			4325: Pixel = 58;
			4326: Pixel = 90;
			4327: Pixel = 85;
			4328: Pixel = 80;
			4329: Pixel = 80;
			4330: Pixel = 147;
			4331: Pixel = 120;
			4332: Pixel = 113;
			4333: Pixel = 114;
			4334: Pixel = 114;
			4335: Pixel = 118;
			4336: Pixel = 127;
			4337: Pixel = 133;
			4338: Pixel = 134;
			4339: Pixel = 119;
			4340: Pixel = 142;
			4341: Pixel = 214;
			4342: Pixel = 207;
			4343: Pixel = 208;
			4344: Pixel = 206;
			4345: Pixel = 203;
			4346: Pixel = 144;
			4347: Pixel = 46;
			4348: Pixel = 43;
			4349: Pixel = 71;
			4350: Pixel = 112;
			4351: Pixel = 78;
			4352: Pixel = 60;
			4353: Pixel = 54;
			4354: Pixel = 94;
			4355: Pixel = 159;
			4356: Pixel = 170;
			4357: Pixel = 173;
			4358: Pixel = 175;
			4359: Pixel = 104;
			4360: Pixel = 100;
			4361: Pixel = 59;
			4362: Pixel = 41;
			4363: Pixel = 74;
			4364: Pixel = 48;
			4365: Pixel = 91;
			4366: Pixel = 59;
			4367: Pixel = 88;
			4368: Pixel = 109;
			4369: Pixel = 117;
			4370: Pixel = 96;
			4371: Pixel = 102;
			4372: Pixel = 110;
			4373: Pixel = 128;
			4374: Pixel = 105;
			4375: Pixel = 66;
			4376: Pixel = 58;
			4377: Pixel = 56;
			4378: Pixel = 56;
			4379: Pixel = 48;
			4380: Pixel = 53;
			4381: Pixel = 50;
			4382: Pixel = 58;
			4383: Pixel = 58;
			4384: Pixel = 58;
			4385: Pixel = 103;
			4386: Pixel = 123;
			4387: Pixel = 124;
			4388: Pixel = 130;
			4389: Pixel = 137;
			4390: Pixel = 140;
			4391: Pixel = 140;
			4392: Pixel = 141;
			4393: Pixel = 159;
			4394: Pixel = 184;
			4395: Pixel = 198;
			4396: Pixel = 209;
			4397: Pixel = 206;
			4398: Pixel = 162;
			4399: Pixel = 66;
			4400: Pixel = 39;
			4401: Pixel = 89;
			4402: Pixel = 79;
			4403: Pixel = 73;
			4404: Pixel = 82;
			4405: Pixel = 146;
			4406: Pixel = 136;
			4407: Pixel = 137;
			4408: Pixel = 127;
			4409: Pixel = 118;
			4410: Pixel = 107;
			4411: Pixel = 100;
			4412: Pixel = 98;
			4413: Pixel = 105;
			4414: Pixel = 101;
			4415: Pixel = 124;
			4416: Pixel = 209;
			4417: Pixel = 204;
			4418: Pixel = 207;
			4419: Pixel = 209;
			4420: Pixel = 142;
			4421: Pixel = 55;
			4422: Pixel = 60;
			4423: Pixel = 81;
			4424: Pixel = 88;
			4425: Pixel = 141;
			4426: Pixel = 134;
			4427: Pixel = 99;
			4428: Pixel = 54;
			4429: Pixel = 85;
			4430: Pixel = 160;
			4431: Pixel = 170;
			4432: Pixel = 174;
			4433: Pixel = 158;
			4434: Pixel = 142;
			4435: Pixel = 106;
			4436: Pixel = 39;
			4437: Pixel = 41;
			4438: Pixel = 85;
			4439: Pixel = 84;
			4440: Pixel = 87;
			4441: Pixel = 72;
			4442: Pixel = 70;
			4443: Pixel = 97;
			4444: Pixel = 82;
			4445: Pixel = 81;
			4446: Pixel = 115;
			4447: Pixel = 139;
			4448: Pixel = 108;
			4449: Pixel = 86;
			4450: Pixel = 96;
			4451: Pixel = 51;
			4452: Pixel = 57;
			4453: Pixel = 59;
			4454: Pixel = 49;
			4455: Pixel = 58;
			4456: Pixel = 53;
			4457: Pixel = 59;
			4458: Pixel = 69;
			4459: Pixel = 57;
			4460: Pixel = 99;
			4461: Pixel = 121;
			4462: Pixel = 124;
			4463: Pixel = 130;
			4464: Pixel = 140;
			4465: Pixel = 139;
			4466: Pixel = 138;
			4467: Pixel = 150;
			4468: Pixel = 165;
			4469: Pixel = 182;
			4470: Pixel = 188;
			4471: Pixel = 191;
			4472: Pixel = 199;
			4473: Pixel = 216;
			4474: Pixel = 206;
			4475: Pixel = 94;
			4476: Pixel = 60;
			4477: Pixel = 75;
			4478: Pixel = 68;
			4479: Pixel = 81;
			4480: Pixel = 149;
			4481: Pixel = 146;
			4482: Pixel = 144;
			4483: Pixel = 140;
			4484: Pixel = 137;
			4485: Pixel = 129;
			4486: Pixel = 119;
			4487: Pixel = 103;
			4488: Pixel = 111;
			4489: Pixel = 108;
			4490: Pixel = 123;
			4491: Pixel = 213;
			4492: Pixel = 209;
			4493: Pixel = 213;
			4494: Pixel = 142;
			4495: Pixel = 53;
			4496: Pixel = 77;
			4497: Pixel = 85;
			4498: Pixel = 93;
			4499: Pixel = 85;
			4500: Pixel = 124;
			4501: Pixel = 151;
			4502: Pixel = 142;
			4503: Pixel = 69;
			4504: Pixel = 83;
			4505: Pixel = 162;
			4506: Pixel = 175;
			4507: Pixel = 175;
			4508: Pixel = 162;
			4509: Pixel = 164;
			4510: Pixel = 74;
			4511: Pixel = 42;
			4512: Pixel = 54;
			4513: Pixel = 60;
			4514: Pixel = 65;
			4515: Pixel = 63;
			4516: Pixel = 63;
			4517: Pixel = 60;
			4518: Pixel = 79;
			4519: Pixel = 64;
			4520: Pixel = 76;
			4521: Pixel = 101;
			4522: Pixel = 139;
			4523: Pixel = 116;
			4524: Pixel = 110;
			4525: Pixel = 113;
			4526: Pixel = 57;
			4527: Pixel = 55;
			4528: Pixel = 62;
			4529: Pixel = 51;
			4530: Pixel = 60;
			4531: Pixel = 55;
			4532: Pixel = 63;
			4533: Pixel = 92;
			4534: Pixel = 60;
			4535: Pixel = 98;
			4536: Pixel = 122;
			4537: Pixel = 125;
			4538: Pixel = 138;
			4539: Pixel = 139;
			4540: Pixel = 139;
			4541: Pixel = 143;
			4542: Pixel = 156;
			4543: Pixel = 164;
			4544: Pixel = 172;
			4545: Pixel = 180;
			4546: Pixel = 186;
			4547: Pixel = 195;
			4548: Pixel = 200;
			4549: Pixel = 214;
			4550: Pixel = 217;
			4551: Pixel = 93;
			4552: Pixel = 49;
			4553: Pixel = 65;
			4554: Pixel = 85;
			4555: Pixel = 150;
			4556: Pixel = 146;
			4557: Pixel = 145;
			4558: Pixel = 142;
			4559: Pixel = 140;
			4560: Pixel = 137;
			4561: Pixel = 131;
			4562: Pixel = 124;
			4563: Pixel = 127;
			4564: Pixel = 119;
			4565: Pixel = 167;
			4566: Pixel = 217;
			4567: Pixel = 212;
			4568: Pixel = 194;
			4569: Pixel = 83;
			4570: Pixel = 76;
			4571: Pixel = 94;
			4572: Pixel = 102;
			4573: Pixel = 100;
			4574: Pixel = 91;
			4575: Pixel = 68;
			4576: Pixel = 144;
			4577: Pixel = 169;
			4578: Pixel = 88;
			4579: Pixel = 78;
			4580: Pixel = 165;
			4581: Pixel = 177;
			4582: Pixel = 177;
			4583: Pixel = 164;
			4584: Pixel = 139;
			4585: Pixel = 59;
			4586: Pixel = 38;
			4587: Pixel = 59;
			4588: Pixel = 55;
			4589: Pixel = 45;
			4590: Pixel = 84;
			4591: Pixel = 53;
			4592: Pixel = 55;
			4593: Pixel = 69;
			4594: Pixel = 78;
			4595: Pixel = 79;
			4596: Pixel = 90;
			4597: Pixel = 112;
			4598: Pixel = 145;
			4599: Pixel = 97;
			4600: Pixel = 111;
			4601: Pixel = 87;
			4602: Pixel = 43;
			4603: Pixel = 63;
			4604: Pixel = 46;
			4605: Pixel = 59;
			4606: Pixel = 54;
			4607: Pixel = 56;
			4608: Pixel = 111;
			4609: Pixel = 67;
			4610: Pixel = 87;
			4611: Pixel = 128;
			4612: Pixel = 133;
			4613: Pixel = 136;
			4614: Pixel = 140;
			4615: Pixel = 140;
			4616: Pixel = 145;
			4617: Pixel = 153;
			4618: Pixel = 160;
			4619: Pixel = 167;
			4620: Pixel = 174;
			4621: Pixel = 182;
			4622: Pixel = 191;
			4623: Pixel = 200;
			4624: Pixel = 204;
			4625: Pixel = 221;
			4626: Pixel = 199;
			4627: Pixel = 56;
			4628: Pixel = 45;
			4629: Pixel = 92;
			4630: Pixel = 149;
			4631: Pixel = 145;
			4632: Pixel = 144;
			4633: Pixel = 142;
			4634: Pixel = 141;
			4635: Pixel = 138;
			4636: Pixel = 134;
			4637: Pixel = 127;
			4638: Pixel = 128;
			4639: Pixel = 139;
			4640: Pixel = 193;
			4641: Pixel = 216;
			4642: Pixel = 215;
			4643: Pixel = 150;
			4644: Pixel = 77;
			4645: Pixel = 95;
			4646: Pixel = 102;
			4647: Pixel = 106;
			4648: Pixel = 94;
			4649: Pixel = 102;
			4650: Pixel = 38;
			4651: Pixel = 129;
			4652: Pixel = 181;
			4653: Pixel = 92;
			4654: Pixel = 69;
			4655: Pixel = 165;
			4656: Pixel = 177;
			4657: Pixel = 178;
			4658: Pixel = 165;
			4659: Pixel = 133;
			4660: Pixel = 63;
			4661: Pixel = 44;
			4662: Pixel = 56;
			4663: Pixel = 45;
			4664: Pixel = 53;
			4665: Pixel = 91;
			4666: Pixel = 55;
			4667: Pixel = 48;
			4668: Pixel = 69;
			4669: Pixel = 67;
			4670: Pixel = 97;
			4671: Pixel = 90;
			4672: Pixel = 97;
			4673: Pixel = 152;
			4674: Pixel = 72;
			4675: Pixel = 107;
			4676: Pixel = 99;
			4677: Pixel = 42;
			4678: Pixel = 71;
			4679: Pixel = 47;
			4680: Pixel = 58;
			4681: Pixel = 49;
			4682: Pixel = 63;
			4683: Pixel = 110;
			4684: Pixel = 70;
			4685: Pixel = 89;
			4686: Pixel = 131;
			4687: Pixel = 131;
			4688: Pixel = 136;
			4689: Pixel = 138;
			4690: Pixel = 141;
			4691: Pixel = 146;
			4692: Pixel = 149;
			4693: Pixel = 156;
			4694: Pixel = 163;
			4695: Pixel = 172;
			4696: Pixel = 180;
			4697: Pixel = 188;
			4698: Pixel = 198;
			4699: Pixel = 207;
			4700: Pixel = 208;
			4701: Pixel = 233;
			4702: Pixel = 127;
			4703: Pixel = 20;
			4704: Pixel = 103;
			4705: Pixel = 152;
			4706: Pixel = 146;
			4707: Pixel = 145;
			4708: Pixel = 142;
			4709: Pixel = 138;
			4710: Pixel = 136;
			4711: Pixel = 133;
			4712: Pixel = 121;
			4713: Pixel = 145;
			4714: Pixel = 189;
			4715: Pixel = 210;
			4716: Pixel = 216;
			4717: Pixel = 204;
			4718: Pixel = 113;
			4719: Pixel = 87;
			4720: Pixel = 102;
			4721: Pixel = 111;
			4722: Pixel = 91;
			4723: Pixel = 97;
			4724: Pixel = 103;
			4725: Pixel = 32;
			4726: Pixel = 115;
			4727: Pixel = 182;
			4728: Pixel = 91;
			4729: Pixel = 66;
			4730: Pixel = 166;
			4731: Pixel = 179;
			4732: Pixel = 180;
			4733: Pixel = 169;
			4734: Pixel = 129;
			4735: Pixel = 54;
			4736: Pixel = 51;
			4737: Pixel = 47;
			4738: Pixel = 38;
			4739: Pixel = 77;
			4740: Pixel = 94;
			4741: Pixel = 42;
			4742: Pixel = 59;
			4743: Pixel = 47;
			4744: Pixel = 51;
			4745: Pixel = 82;
			4746: Pixel = 94;
			4747: Pixel = 87;
			4748: Pixel = 148;
			4749: Pixel = 107;
			4750: Pixel = 121;
			4751: Pixel = 92;
			4752: Pixel = 49;
			4753: Pixel = 65;
			4754: Pixel = 52;
			4755: Pixel = 54;
			4756: Pixel = 50;
			4757: Pixel = 81;
			4758: Pixel = 124;
			4759: Pixel = 79;
			4760: Pixel = 94;
			4761: Pixel = 133;
			4762: Pixel = 135;
			4763: Pixel = 137;
			4764: Pixel = 136;
			4765: Pixel = 138;
			4766: Pixel = 144;
			4767: Pixel = 147;
			4768: Pixel = 154;
			4769: Pixel = 161;
			4770: Pixel = 168;
			4771: Pixel = 177;
			4772: Pixel = 186;
			4773: Pixel = 196;
			4774: Pixel = 206;
			4775: Pixel = 209;
			4776: Pixel = 222;
			4777: Pixel = 194;
			4778: Pixel = 29;
			4779: Pixel = 109;
			4780: Pixel = 154;
			4781: Pixel = 145;
			4782: Pixel = 145;
			4783: Pixel = 141;
			4784: Pixel = 137;
			4785: Pixel = 132;
			4786: Pixel = 126;
			4787: Pixel = 125;
			4788: Pixel = 197;
			4789: Pixel = 212;
			4790: Pixel = 212;
			4791: Pixel = 219;
			4792: Pixel = 167;
			4793: Pixel = 91;
			4794: Pixel = 93;
			4795: Pixel = 112;
			4796: Pixel = 102;
			4797: Pixel = 93;
			4798: Pixel = 104;
			4799: Pixel = 100;
			4800: Pixel = 27;
			4801: Pixel = 107;
			4802: Pixel = 182;
			4803: Pixel = 103;
			4804: Pixel = 64;
			4805: Pixel = 165;
			4806: Pixel = 177;
			4807: Pixel = 176;
			4808: Pixel = 167;
			4809: Pixel = 120;
			4810: Pixel = 55;
			4811: Pixel = 45;
			4812: Pixel = 46;
			4813: Pixel = 53;
			4814: Pixel = 76;
			4815: Pixel = 76;
			4816: Pixel = 48;
			4817: Pixel = 57;
			4818: Pixel = 45;
			4819: Pixel = 56;
			4820: Pixel = 62;
			4821: Pixel = 82;
			4822: Pixel = 123;
			4823: Pixel = 126;
			4824: Pixel = 115;
			4825: Pixel = 141;
			4826: Pixel = 85;
			4827: Pixel = 68;
			4828: Pixel = 63;
			4829: Pixel = 57;
			4830: Pixel = 51;
			4831: Pixel = 58;
			4832: Pixel = 108;
			4833: Pixel = 130;
			4834: Pixel = 76;
			4835: Pixel = 101;
			4836: Pixel = 133;
			4837: Pixel = 136;
			4838: Pixel = 139;
			4839: Pixel = 136;
			4840: Pixel = 137;
			4841: Pixel = 141;
			4842: Pixel = 145;
			4843: Pixel = 152;
			4844: Pixel = 158;
			4845: Pixel = 165;
			4846: Pixel = 174;
			4847: Pixel = 185;
			4848: Pixel = 194;
			4849: Pixel = 204;
			4850: Pixel = 209;
			4851: Pixel = 212;
			4852: Pixel = 223;
			4853: Pixel = 70;
			4854: Pixel = 109;
			4855: Pixel = 154;
			4856: Pixel = 143;
			4857: Pixel = 141;
			4858: Pixel = 139;
			4859: Pixel = 138;
			4860: Pixel = 133;
			4861: Pixel = 122;
			4862: Pixel = 138;
			4863: Pixel = 212;
			4864: Pixel = 209;
			4865: Pixel = 216;
			4866: Pixel = 206;
			4867: Pixel = 133;
			4868: Pixel = 97;
			4869: Pixel = 99;
			4870: Pixel = 112;
			4871: Pixel = 94;
			4872: Pixel = 100;
			4873: Pixel = 101;
			4874: Pixel = 88;
			4875: Pixel = 27;
			4876: Pixel = 97;
			4877: Pixel = 182;
			4878: Pixel = 112;
			4879: Pixel = 64;
			4880: Pixel = 162;
			4881: Pixel = 177;
			4882: Pixel = 176;
			4883: Pixel = 168;
			4884: Pixel = 126;
			4885: Pixel = 52;
			4886: Pixel = 45;
			4887: Pixel = 46;
			4888: Pixel = 56;
			4889: Pixel = 53;
			4890: Pixel = 69;
			4891: Pixel = 51;
			4892: Pixel = 54;
			4893: Pixel = 45;
			4894: Pixel = 61;
			4895: Pixel = 67;
			4896: Pixel = 63;
			4897: Pixel = 120;
			4898: Pixel = 119;
			4899: Pixel = 82;
			4900: Pixel = 57;
			4901: Pixel = 68;
			4902: Pixel = 83;
			4903: Pixel = 89;
			4904: Pixel = 63;
			4905: Pixel = 47;
			4906: Pixel = 76;
			4907: Pixel = 120;
			4908: Pixel = 127;
			4909: Pixel = 76;
			4910: Pixel = 113;
			4911: Pixel = 135;
			4912: Pixel = 137;
			4913: Pixel = 140;
			4914: Pixel = 136;
			4915: Pixel = 134;
			4916: Pixel = 139;
			4917: Pixel = 143;
			4918: Pixel = 149;
			4919: Pixel = 156;
			4920: Pixel = 162;
			4921: Pixel = 170;
			4922: Pixel = 181;
			4923: Pixel = 192;
			4924: Pixel = 201;
			4925: Pixel = 207;
			4926: Pixel = 209;
			4927: Pixel = 227;
			4928: Pixel = 123;
			4929: Pixel = 112;
			4930: Pixel = 155;
			4931: Pixel = 144;
			4932: Pixel = 140;
			4933: Pixel = 138;
			4934: Pixel = 138;
			4935: Pixel = 133;
			4936: Pixel = 123;
			4937: Pixel = 145;
			4938: Pixel = 211;
			4939: Pixel = 205;
			4940: Pixel = 219;
			4941: Pixel = 176;
			4942: Pixel = 115;
			4943: Pixel = 103;
			4944: Pixel = 100;
			4945: Pixel = 98;
			4946: Pixel = 91;
			4947: Pixel = 103;
			4948: Pixel = 93;
			4949: Pixel = 90;
			4950: Pixel = 30;
			4951: Pixel = 82;
			4952: Pixel = 175;
			4953: Pixel = 121;
			4954: Pixel = 71;
			4955: Pixel = 158;
			4956: Pixel = 178;
			4957: Pixel = 178;
			4958: Pixel = 168;
			4959: Pixel = 133;
			4960: Pixel = 58;
			4961: Pixel = 42;
			4962: Pixel = 60;
			4963: Pixel = 58;
			4964: Pixel = 50;
			4965: Pixel = 60;
			4966: Pixel = 53;
			4967: Pixel = 58;
			4968: Pixel = 51;
			4969: Pixel = 62;
			4970: Pixel = 69;
			4971: Pixel = 77;
			4972: Pixel = 115;
			4973: Pixel = 99;
			4974: Pixel = 105;
			4975: Pixel = 98;
			4976: Pixel = 47;
			4977: Pixel = 51;
			4978: Pixel = 55;
			4979: Pixel = 51;
			4980: Pixel = 52;
			4981: Pixel = 95;
			4982: Pixel = 125;
			4983: Pixel = 114;
			4984: Pixel = 77;
			4985: Pixel = 127;
			4986: Pixel = 139;
			4987: Pixel = 140;
			4988: Pixel = 140;
			4989: Pixel = 137;
			4990: Pixel = 136;
			4991: Pixel = 137;
			4992: Pixel = 142;
			4993: Pixel = 147;
			4994: Pixel = 153;
			4995: Pixel = 159;
			4996: Pixel = 165;
			4997: Pixel = 176;
			4998: Pixel = 189;
			4999: Pixel = 198;
			5000: Pixel = 205;
			5001: Pixel = 208;
			5002: Pixel = 220;
			5003: Pixel = 177;
			5004: Pixel = 126;
			5005: Pixel = 141;
			5006: Pixel = 142;
			5007: Pixel = 146;
			5008: Pixel = 144;
			5009: Pixel = 141;
			5010: Pixel = 134;
			5011: Pixel = 133;
			5012: Pixel = 140;
			5013: Pixel = 162;
			5014: Pixel = 199;
			5015: Pixel = 219;
			5016: Pixel = 155;
			5017: Pixel = 106;
			5018: Pixel = 98;
			5019: Pixel = 95;
			5020: Pixel = 82;
			5021: Pixel = 103;
			5022: Pixel = 93;
			5023: Pixel = 93;
			5024: Pixel = 94;
			5025: Pixel = 31;
			5026: Pixel = 73;
			5027: Pixel = 171;
			5028: Pixel = 131;
			5029: Pixel = 74;
			5030: Pixel = 154;
			5031: Pixel = 176;
			5032: Pixel = 177;
			5033: Pixel = 168;
			5034: Pixel = 132;
			5035: Pixel = 68;
			5036: Pixel = 45;
			5037: Pixel = 55;
			5038: Pixel = 45;
			5039: Pixel = 57;
			5040: Pixel = 60;
			5041: Pixel = 61;
			5042: Pixel = 50;
			5043: Pixel = 50;
			5044: Pixel = 58;
			5045: Pixel = 78;
			5046: Pixel = 87;
			5047: Pixel = 55;
			5048: Pixel = 75;
			5049: Pixel = 86;
			5050: Pixel = 116;
			5051: Pixel = 47;
			5052: Pixel = 50;
			5053: Pixel = 47;
			5054: Pixel = 43;
			5055: Pixel = 68;
			5056: Pixel = 108;
			5057: Pixel = 129;
			5058: Pixel = 89;
			5059: Pixel = 89;
			5060: Pixel = 137;
			5061: Pixel = 137;
			5062: Pixel = 142;
			5063: Pixel = 142;
			5064: Pixel = 140;
			5065: Pixel = 137;
			5066: Pixel = 137;
			5067: Pixel = 141;
			5068: Pixel = 147;
			5069: Pixel = 150;
			5070: Pixel = 155;
			5071: Pixel = 163;
			5072: Pixel = 172;
			5073: Pixel = 184;
			5074: Pixel = 194;
			5075: Pixel = 203;
			5076: Pixel = 210;
			5077: Pixel = 213;
			5078: Pixel = 213;
			5079: Pixel = 122;
			5080: Pixel = 83;
			5081: Pixel = 102;
			5082: Pixel = 120;
			5083: Pixel = 134;
			5084: Pixel = 140;
			5085: Pixel = 142;
			5086: Pixel = 151;
			5087: Pixel = 140;
			5088: Pixel = 133;
			5089: Pixel = 204;
			5090: Pixel = 211;
			5091: Pixel = 134;
			5092: Pixel = 92;
			5093: Pixel = 94;
			5094: Pixel = 82;
			5095: Pixel = 93;
			5096: Pixel = 99;
			5097: Pixel = 92;
			5098: Pixel = 97;
			5099: Pixel = 76;
			5100: Pixel = 27;
			5101: Pixel = 62;
			5102: Pixel = 174;
			5103: Pixel = 146;
			5104: Pixel = 74;
			5105: Pixel = 148;
			5106: Pixel = 175;
			5107: Pixel = 177;
			5108: Pixel = 170;
			5109: Pixel = 120;
			5110: Pixel = 73;
			5111: Pixel = 45;
			5112: Pixel = 44;
			5113: Pixel = 55;
			5114: Pixel = 57;
			5115: Pixel = 55;
			5116: Pixel = 63;
			5117: Pixel = 48;
			5118: Pixel = 48;
			5119: Pixel = 52;
			5120: Pixel = 76;
			5121: Pixel = 127;
			5122: Pixel = 83;
			5123: Pixel = 77;
			5124: Pixel = 76;
			5125: Pixel = 54;
			5126: Pixel = 46;
			5127: Pixel = 46;
			5128: Pixel = 41;
			5129: Pixel = 53;
			5130: Pixel = 92;
			5131: Pixel = 121;
			5132: Pixel = 112;
			5133: Pixel = 62;
			5134: Pixel = 119;
			5135: Pixel = 136;
			5136: Pixel = 137;
			5137: Pixel = 142;
			5138: Pixel = 141;
			5139: Pixel = 141;
			5140: Pixel = 138;
			5141: Pixel = 135;
			5142: Pixel = 138;
			5143: Pixel = 143;
			5144: Pixel = 148;
			5145: Pixel = 153;
			5146: Pixel = 160;
			5147: Pixel = 168;
			5148: Pixel = 178;
			5149: Pixel = 190;
			5150: Pixel = 201;
			5151: Pixel = 208;
			5152: Pixel = 210;
			5153: Pixel = 224;
			5154: Pixel = 124;
			5155: Pixel = 75;
			5156: Pixel = 81;
			5157: Pixel = 76;
			5158: Pixel = 77;
			5159: Pixel = 82;
			5160: Pixel = 102;
			5161: Pixel = 140;
			5162: Pixel = 153;
			5163: Pixel = 159;
			5164: Pixel = 218;
			5165: Pixel = 182;
			5166: Pixel = 91;
			5167: Pixel = 74;
			5168: Pixel = 85;
			5169: Pixel = 88;
			5170: Pixel = 100;
			5171: Pixel = 90;
			5172: Pixel = 100;
			5173: Pixel = 91;
			5174: Pixel = 58;
			5175: Pixel = 59;
			5176: Pixel = 76;
			5177: Pixel = 170;
			5178: Pixel = 163;
			5179: Pixel = 82;
			5180: Pixel = 146;
			5181: Pixel = 175;
			5182: Pixel = 178;
			5183: Pixel = 170;
			5184: Pixel = 115;
			5185: Pixel = 66;
			5186: Pixel = 45;
			5187: Pixel = 52;
			5188: Pixel = 53;
			5189: Pixel = 51;
			5190: Pixel = 57;
			5191: Pixel = 62;
			5192: Pixel = 55;
			5193: Pixel = 46;
			5194: Pixel = 50;
			5195: Pixel = 47;
			5196: Pixel = 86;
			5197: Pixel = 138;
			5198: Pixel = 110;
			5199: Pixel = 73;
			5200: Pixel = 41;
			5201: Pixel = 47;
			5202: Pixel = 41;
			5203: Pixel = 41;
			5204: Pixel = 71;
			5205: Pixel = 112;
			5206: Pixel = 124;
			5207: Pixel = 63;
			5208: Pixel = 87;
			5209: Pixel = 137;
			5210: Pixel = 136;
			5211: Pixel = 138;
			5212: Pixel = 139;
			5213: Pixel = 142;
			5214: Pixel = 143;
			5215: Pixel = 140;
			5216: Pixel = 137;
			5217: Pixel = 137;
			5218: Pixel = 139;
			5219: Pixel = 145;
			5220: Pixel = 151;
			5221: Pixel = 156;
			5222: Pixel = 163;
			5223: Pixel = 175;
			5224: Pixel = 186;
			5225: Pixel = 198;
			5226: Pixel = 205;
			5227: Pixel = 208;
			5228: Pixel = 223;
			5229: Pixel = 164;
			5230: Pixel = 90;
			5231: Pixel = 106;
			5232: Pixel = 91;
			5233: Pixel = 72;
			5234: Pixel = 50;
			5235: Pixel = 31;
			5236: Pixel = 116;
			5237: Pixel = 192;
			5238: Pixel = 179;
			5239: Pixel = 220;
			5240: Pixel = 122;
			5241: Pixel = 58;
			5242: Pixel = 74;
			5243: Pixel = 82;
			5244: Pixel = 104;
			5245: Pixel = 85;
			5246: Pixel = 88;
			5247: Pixel = 105;
			5248: Pixel = 79;
			5249: Pixel = 55;
			5250: Pixel = 92;
			5251: Pixel = 108;
			5252: Pixel = 167;
			5253: Pixel = 172;
			5254: Pixel = 95;
			5255: Pixel = 143;
			5256: Pixel = 177;
			5257: Pixel = 181;
			5258: Pixel = 168;
			5259: Pixel = 115;
			5260: Pixel = 63;
			5261: Pixel = 46;
			5262: Pixel = 50;
			5263: Pixel = 49;
			5264: Pixel = 50;
			5265: Pixel = 52;
			5266: Pixel = 62;
			5267: Pixel = 58;
			5268: Pixel = 45;
			5269: Pixel = 59;
			5270: Pixel = 61;
			5271: Pixel = 55;
			5272: Pixel = 96;
			5273: Pixel = 113;
			5274: Pixel = 71;
			5275: Pixel = 43;
			5276: Pixel = 42;
			5277: Pixel = 39;
			5278: Pixel = 62;
			5279: Pixel = 100;
			5280: Pixel = 113;
			5281: Pixel = 66;
			5282: Pixel = 72;
			5283: Pixel = 128;
			5284: Pixel = 133;
			5285: Pixel = 137;
			5286: Pixel = 139;
			5287: Pixel = 139;
			5288: Pixel = 141;
			5289: Pixel = 142;
			5290: Pixel = 141;
			5291: Pixel = 139;
			5292: Pixel = 138;
			5293: Pixel = 139;
			5294: Pixel = 141;
			5295: Pixel = 147;
			5296: Pixel = 153;
			5297: Pixel = 161;
			5298: Pixel = 168;
			5299: Pixel = 180;
			5300: Pixel = 193;
			5301: Pixel = 202;
			5302: Pixel = 208;
			5303: Pixel = 216;
			5304: Pixel = 196;
			5305: Pixel = 93;
			5306: Pixel = 107;
			5307: Pixel = 103;
			5308: Pixel = 91;
			5309: Pixel = 76;
			5310: Pixel = 45;
			5311: Pixel = 121;
			5312: Pixel = 206;
			5313: Pixel = 192;
			5314: Pixel = 143;
			5315: Pixel = 54;
			5316: Pixel = 64;
			5317: Pixel = 74;
			5318: Pixel = 101;
			5319: Pixel = 87;
			5320: Pixel = 75;
			5321: Pixel = 101;
			5322: Pixel = 104;
			5323: Pixel = 76;
			5324: Pixel = 63;
			5325: Pixel = 80;
			5326: Pixel = 111;
			5327: Pixel = 159;
			5328: Pixel = 171;
			5329: Pixel = 101;
			5330: Pixel = 141;
			5331: Pixel = 177;
			5332: Pixel = 182;
			5333: Pixel = 170;
			5334: Pixel = 107;
			5335: Pixel = 52;
			5336: Pixel = 47;
			5337: Pixel = 53;
			5338: Pixel = 54;
			5339: Pixel = 51;
			5340: Pixel = 58;
			5341: Pixel = 70;
			5342: Pixel = 79;
			5343: Pixel = 58;
			5344: Pixel = 62;
			5345: Pixel = 66;
			5346: Pixel = 69;
			5347: Pixel = 93;
			5348: Pixel = 99;
			5349: Pixel = 51;
			5350: Pixel = 43;
			5351: Pixel = 43;
			5352: Pixel = 45;
			5353: Pixel = 69;
			5354: Pixel = 73;
			5355: Pixel = 64;
			5356: Pixel = 86;
			5357: Pixel = 122;
			5358: Pixel = 128;
			5359: Pixel = 133;
			5360: Pixel = 136;
			5361: Pixel = 138;
			5362: Pixel = 139;
			5363: Pixel = 141;
			5364: Pixel = 143;
			5365: Pixel = 145;
			5366: Pixel = 143;
			5367: Pixel = 140;
			5368: Pixel = 139;
			5369: Pixel = 140;
			5370: Pixel = 144;
			5371: Pixel = 150;
			5372: Pixel = 158;
			5373: Pixel = 166;
			5374: Pixel = 174;
			5375: Pixel = 186;
			5376: Pixel = 198;
			5377: Pixel = 206;
			5378: Pixel = 211;
			5379: Pixel = 216;
			5380: Pixel = 111;
			5381: Pixel = 93;
			5382: Pixel = 104;
			5383: Pixel = 99;
			5384: Pixel = 93;
			5385: Pixel = 87;
			5386: Pixel = 126;
			5387: Pixel = 199;
			5388: Pixel = 122;
			5389: Pixel = 63;
			5390: Pixel = 67;
			5391: Pixel = 74;
			5392: Pixel = 101;
			5393: Pixel = 94;
			5394: Pixel = 67;
			5395: Pixel = 89;
			5396: Pixel = 113;
			5397: Pixel = 94;
			5398: Pixel = 68;
			5399: Pixel = 65;
			5400: Pixel = 57;
			5401: Pixel = 82;
			5402: Pixel = 146;
			5403: Pixel = 174;
			5404: Pixel = 110;
			5405: Pixel = 138;
			5406: Pixel = 178;
			5407: Pixel = 182;
			5408: Pixel = 176;
			5409: Pixel = 89;
			5410: Pixel = 45;
			5411: Pixel = 48;
			5412: Pixel = 56;
			5413: Pixel = 59;
			5414: Pixel = 59;
			5415: Pixel = 58;
			5416: Pixel = 61;
			5417: Pixel = 86;
			5418: Pixel = 83;
			5419: Pixel = 66;
			5420: Pixel = 67;
			5421: Pixel = 72;
			5422: Pixel = 90;
			5423: Pixel = 112;
			5424: Pixel = 52;
			5425: Pixel = 45;
			5426: Pixel = 43;
			5427: Pixel = 50;
			5428: Pixel = 70;
			5429: Pixel = 86;
			5430: Pixel = 112;
			5431: Pixel = 126;
			5432: Pixel = 127;
			5433: Pixel = 127;
			5434: Pixel = 130;
			5435: Pixel = 135;
			5436: Pixel = 136;
			5437: Pixel = 139;
			5438: Pixel = 141;
			5439: Pixel = 143;
			5440: Pixel = 146;
			5441: Pixel = 144;
			5442: Pixel = 143;
			5443: Pixel = 141;
			5444: Pixel = 141;
			5445: Pixel = 144;
			5446: Pixel = 149;
			5447: Pixel = 155;
			5448: Pixel = 162;
			5449: Pixel = 173;
			5450: Pixel = 183;
			5451: Pixel = 192;
			5452: Pixel = 201;
			5453: Pixel = 208;
			5454: Pixel = 222;
			5455: Pixel = 141;
			5456: Pixel = 79;
			5457: Pixel = 105;
			5458: Pixel = 108;
			5459: Pixel = 108;
			5460: Pixel = 113;
			5461: Pixel = 114;
			5462: Pixel = 110;
			5463: Pixel = 83;
			5464: Pixel = 89;
			5465: Pixel = 77;
			5466: Pixel = 92;
			5467: Pixel = 97;
			5468: Pixel = 69;
			5469: Pixel = 72;
			5470: Pixel = 112;
			5471: Pixel = 114;
			5472: Pixel = 82;
			5473: Pixel = 60;
			5474: Pixel = 54;
			5475: Pixel = 54;
			5476: Pixel = 59;
			5477: Pixel = 151;
			5478: Pixel = 206;
			5479: Pixel = 135;
			5480: Pixel = 136;
			5481: Pixel = 178;
			5482: Pixel = 184;
			5483: Pixel = 167;
			5484: Pixel = 75;
			5485: Pixel = 49;
			5486: Pixel = 49;
			5487: Pixel = 56;
			5488: Pixel = 61;
			5489: Pixel = 60;
			5490: Pixel = 66;
			5491: Pixel = 64;
			5492: Pixel = 73;
			5493: Pixel = 102;
			5494: Pixel = 69;
			5495: Pixel = 73;
			5496: Pixel = 65;
			5497: Pixel = 76;
			5498: Pixel = 90;
			5499: Pixel = 65;
			5500: Pixel = 38;
			5501: Pixel = 53;
			5502: Pixel = 84;
			5503: Pixel = 110;
			5504: Pixel = 119;
			5505: Pixel = 121;
			5506: Pixel = 125;
			5507: Pixel = 127;
			5508: Pixel = 129;
			5509: Pixel = 130;
			5510: Pixel = 134;
			5511: Pixel = 136;
			5512: Pixel = 138;
			5513: Pixel = 140;
			5514: Pixel = 141;
			5515: Pixel = 144;
			5516: Pixel = 146;
			5517: Pixel = 146;
			5518: Pixel = 146;
			5519: Pixel = 145;
			5520: Pixel = 146;
			5521: Pixel = 149;
			5522: Pixel = 153;
			5523: Pixel = 161;
			5524: Pixel = 168;
			5525: Pixel = 178;
			5526: Pixel = 187;
			5527: Pixel = 197;
			5528: Pixel = 204;
			5529: Pixel = 217;
			5530: Pixel = 173;
			5531: Pixel = 76;
			5532: Pixel = 102;
			5533: Pixel = 110;
			5534: Pixel = 119;
			5535: Pixel = 118;
			5536: Pixel = 111;
			5537: Pixel = 103;
			5538: Pixel = 115;
			5539: Pixel = 100;
			5540: Pixel = 91;
			5541: Pixel = 92;
			5542: Pixel = 72;
			5543: Pixel = 73;
			5544: Pixel = 103;
			5545: Pixel = 123;
			5546: Pixel = 96;
			5547: Pixel = 62;
			5548: Pixel = 54;
			5549: Pixel = 59;
			5550: Pixel = 50;
			5551: Pixel = 49;
			5552: Pixel = 154;
			5553: Pixel = 212;
			5554: Pixel = 148;
			5555: Pixel = 136;
			5556: Pixel = 177;
			5557: Pixel = 183;
			5558: Pixel = 164;
			5559: Pixel = 74;
			5560: Pixel = 44;
			5561: Pixel = 54;
			5562: Pixel = 60;
			5563: Pixel = 70;
			5564: Pixel = 62;
			5565: Pixel = 87;
			5566: Pixel = 66;
			5567: Pixel = 76;
			5568: Pixel = 87;
			5569: Pixel = 84;
			5570: Pixel = 80;
			5571: Pixel = 59;
			5572: Pixel = 67;
			5573: Pixel = 67;
			5574: Pixel = 94;
			5575: Pixel = 59;
			5576: Pixel = 75;
			5577: Pixel = 100;
			5578: Pixel = 113;
			5579: Pixel = 119;
			5580: Pixel = 123;
			5581: Pixel = 126;
			5582: Pixel = 127;
			5583: Pixel = 130;
			5584: Pixel = 131;
			5585: Pixel = 133;
			5586: Pixel = 136;
			5587: Pixel = 135;
			5588: Pixel = 139;
			5589: Pixel = 141;
			5590: Pixel = 145;
			5591: Pixel = 144;
			5592: Pixel = 145;
			5593: Pixel = 148;
			5594: Pixel = 149;
			5595: Pixel = 148;
			5596: Pixel = 152;
			5597: Pixel = 155;
			5598: Pixel = 161;
			5599: Pixel = 166;
			5600: Pixel = 174;
			5601: Pixel = 185;
			5602: Pixel = 194;
			5603: Pixel = 201;
			5604: Pixel = 211;
			5605: Pixel = 200;
			5606: Pixel = 94;
			5607: Pixel = 90;
			5608: Pixel = 105;
			5609: Pixel = 120;
			5610: Pixel = 125;
			5611: Pixel = 118;
			5612: Pixel = 129;
			5613: Pixel = 122;
			5614: Pixel = 94;
			5615: Pixel = 85;
			5616: Pixel = 84;
			5617: Pixel = 82;
			5618: Pixel = 92;
			5619: Pixel = 129;
			5620: Pixel = 111;
			5621: Pixel = 65;
			5622: Pixel = 46;
			5623: Pixel = 63;
			5624: Pixel = 93;
		endcase
	end
endmodule