module InHandle(
	input wire			nReset,                                                      // Common to all
	input wire			Clk,                                                        // Common to all
	output reg	[7:0]	Pixel,
	output reg			Frame,
	output reg			Line
);

	parameter COLS = 100;
	parameter ROWS = 100;
	
	reg [7:0] col;
	reg [7:0] row;
	
	always @ (posedge Clk or negedge nReset) begin
		if(!nReset) begin   
			Frame <= 0;
	    	Line  <= 0;							
			row <= ROWS-1;
			col <= COLS-1;						// Zero on first pixel	
		end else begin
			if(col == (COLS-1)) begin			// Get ready for next column
	    		Line <= 1;
				col <= 0;
				row <= row + 1;
				if(row == (ROWS-1)) begin		// Get ready for next row
					Frame <= 1;
					row <= 0;
				end
			end else begin
				Line <= 0;
				Frame <= 0;
				col = col + 1;
			end
		end
	end

	always @ (*) begin
		case(col + (row*COLS))


			0: Pixel = 161;
			1: Pixel = 161;
			2: Pixel = 159;
			3: Pixel = 157;
			4: Pixel = 156;
			5: Pixel = 154;
			6: Pixel = 155;
			7: Pixel = 162;
			8: Pixel = 170;
			9: Pixel = 172;
			10: Pixel = 165;
			11: Pixel = 142;
			12: Pixel = 103;
			13: Pixel = 94;
			14: Pixel = 103;
			15: Pixel = 106;
			16: Pixel = 107;
			17: Pixel = 108;
			18: Pixel = 109;
			19: Pixel = 106;
			20: Pixel = 109;
			21: Pixel = 117;
			22: Pixel = 121;
			23: Pixel = 125;
			24: Pixel = 128;
			25: Pixel = 130;
			26: Pixel = 131;
			27: Pixel = 131;
			28: Pixel = 129;
			29: Pixel = 129;
			30: Pixel = 131;
			31: Pixel = 132;
			32: Pixel = 133;
			33: Pixel = 133;
			34: Pixel = 134;
			35: Pixel = 132;
			36: Pixel = 133;
			37: Pixel = 133;
			38: Pixel = 135;
			39: Pixel = 134;
			40: Pixel = 135;
			41: Pixel = 133;
			42: Pixel = 130;
			43: Pixel = 130;
			44: Pixel = 132;
			45: Pixel = 131;
			46: Pixel = 131;
			47: Pixel = 134;
			48: Pixel = 133;
			49: Pixel = 133;
			50: Pixel = 135;
			51: Pixel = 129;
			52: Pixel = 131;
			53: Pixel = 129;
			54: Pixel = 131;
			55: Pixel = 129;
			56: Pixel = 130;
			57: Pixel = 128;
			58: Pixel = 127;
			59: Pixel = 124;
			60: Pixel = 120;
			61: Pixel = 112;
			62: Pixel = 105;
			63: Pixel = 127;
			64: Pixel = 146;
			65: Pixel = 157;
			66: Pixel = 159;
			67: Pixel = 151;
			68: Pixel = 152;
			69: Pixel = 154;
			70: Pixel = 156;
			71: Pixel = 153;
			72: Pixel = 153;
			73: Pixel = 152;
			74: Pixel = 153;
			75: Pixel = 155;
			76: Pixel = 157;
			77: Pixel = 155;
			78: Pixel = 162;
			79: Pixel = 206;
			80: Pixel = 216;
			81: Pixel = 218;
			82: Pixel = 149;
			83: Pixel = 98;
			84: Pixel = 115;
			85: Pixel = 121;
			86: Pixel = 120;
			87: Pixel = 122;
			88: Pixel = 122;
			89: Pixel = 121;
			90: Pixel = 122;
			91: Pixel = 124;
			92: Pixel = 124;
			93: Pixel = 122;
			94: Pixel = 125;
			95: Pixel = 125;
			96: Pixel = 123;
			97: Pixel = 112;
			98: Pixel = 145;
			99: Pixel = 163;
			100: Pixel = 158;
			101: Pixel = 158;
			102: Pixel = 156;
			103: Pixel = 155;
			104: Pixel = 154;
			105: Pixel = 153;
			106: Pixel = 153;
			107: Pixel = 162;
			108: Pixel = 170;
			109: Pixel = 172;
			110: Pixel = 162;
			111: Pixel = 136;
			112: Pixel = 102;
			113: Pixel = 90;
			114: Pixel = 99;
			115: Pixel = 104;
			116: Pixel = 103;
			117: Pixel = 105;
			118: Pixel = 104;
			119: Pixel = 105;
			120: Pixel = 109;
			121: Pixel = 116;
			122: Pixel = 122;
			123: Pixel = 124;
			124: Pixel = 125;
			125: Pixel = 129;
			126: Pixel = 129;
			127: Pixel = 130;
			128: Pixel = 130;
			129: Pixel = 130;
			130: Pixel = 130;
			131: Pixel = 132;
			132: Pixel = 134;
			133: Pixel = 133;
			134: Pixel = 133;
			135: Pixel = 131;
			136: Pixel = 131;
			137: Pixel = 132;
			138: Pixel = 132;
			139: Pixel = 131;
			140: Pixel = 131;
			141: Pixel = 132;
			142: Pixel = 129;
			143: Pixel = 129;
			144: Pixel = 132;
			145: Pixel = 128;
			146: Pixel = 130;
			147: Pixel = 132;
			148: Pixel = 131;
			149: Pixel = 130;
			150: Pixel = 132;
			151: Pixel = 129;
			152: Pixel = 128;
			153: Pixel = 128;
			154: Pixel = 127;
			155: Pixel = 127;
			156: Pixel = 129;
			157: Pixel = 128;
			158: Pixel = 126;
			159: Pixel = 124;
			160: Pixel = 119;
			161: Pixel = 112;
			162: Pixel = 104;
			163: Pixel = 119;
			164: Pixel = 141;
			165: Pixel = 153;
			166: Pixel = 159;
			167: Pixel = 154;
			168: Pixel = 152;
			169: Pixel = 154;
			170: Pixel = 154;
			171: Pixel = 155;
			172: Pixel = 153;
			173: Pixel = 153;
			174: Pixel = 153;
			175: Pixel = 154;
			176: Pixel = 155;
			177: Pixel = 154;
			178: Pixel = 152;
			179: Pixel = 192;
			180: Pixel = 215;
			181: Pixel = 220;
			182: Pixel = 181;
			183: Pixel = 105;
			184: Pixel = 110;
			185: Pixel = 119;
			186: Pixel = 120;
			187: Pixel = 121;
			188: Pixel = 121;
			189: Pixel = 120;
			190: Pixel = 123;
			191: Pixel = 123;
			192: Pixel = 123;
			193: Pixel = 123;
			194: Pixel = 125;
			195: Pixel = 125;
			196: Pixel = 125;
			197: Pixel = 127;
			198: Pixel = 108;
			199: Pixel = 72;
			200: Pixel = 156;
			201: Pixel = 155;
			202: Pixel = 155;
			203: Pixel = 156;
			204: Pixel = 154;
			205: Pixel = 153;
			206: Pixel = 157;
			207: Pixel = 166;
			208: Pixel = 169;
			209: Pixel = 169;
			210: Pixel = 159;
			211: Pixel = 133;
			212: Pixel = 100;
			213: Pixel = 89;
			214: Pixel = 98;
			215: Pixel = 103;
			216: Pixel = 106;
			217: Pixel = 105;
			218: Pixel = 103;
			219: Pixel = 102;
			220: Pixel = 109;
			221: Pixel = 115;
			222: Pixel = 120;
			223: Pixel = 123;
			224: Pixel = 125;
			225: Pixel = 127;
			226: Pixel = 128;
			227: Pixel = 130;
			228: Pixel = 131;
			229: Pixel = 129;
			230: Pixel = 129;
			231: Pixel = 131;
			232: Pixel = 131;
			233: Pixel = 133;
			234: Pixel = 132;
			235: Pixel = 131;
			236: Pixel = 132;
			237: Pixel = 131;
			238: Pixel = 131;
			239: Pixel = 130;
			240: Pixel = 131;
			241: Pixel = 131;
			242: Pixel = 130;
			243: Pixel = 129;
			244: Pixel = 130;
			245: Pixel = 129;
			246: Pixel = 130;
			247: Pixel = 133;
			248: Pixel = 132;
			249: Pixel = 130;
			250: Pixel = 130;
			251: Pixel = 130;
			252: Pixel = 129;
			253: Pixel = 128;
			254: Pixel = 127;
			255: Pixel = 127;
			256: Pixel = 127;
			257: Pixel = 128;
			258: Pixel = 128;
			259: Pixel = 125;
			260: Pixel = 120;
			261: Pixel = 114;
			262: Pixel = 108;
			263: Pixel = 106;
			264: Pixel = 131;
			265: Pixel = 149;
			266: Pixel = 158;
			267: Pixel = 159;
			268: Pixel = 156;
			269: Pixel = 158;
			270: Pixel = 159;
			271: Pixel = 158;
			272: Pixel = 155;
			273: Pixel = 155;
			274: Pixel = 154;
			275: Pixel = 153;
			276: Pixel = 152;
			277: Pixel = 153;
			278: Pixel = 149;
			279: Pixel = 162;
			280: Pixel = 207;
			281: Pixel = 217;
			282: Pixel = 218;
			283: Pixel = 146;
			284: Pixel = 101;
			285: Pixel = 115;
			286: Pixel = 118;
			287: Pixel = 120;
			288: Pixel = 121;
			289: Pixel = 119;
			290: Pixel = 121;
			291: Pixel = 121;
			292: Pixel = 122;
			293: Pixel = 123;
			294: Pixel = 124;
			295: Pixel = 126;
			296: Pixel = 135;
			297: Pixel = 101;
			298: Pixel = 48;
			299: Pixel = 41;
			300: Pixel = 156;
			301: Pixel = 156;
			302: Pixel = 156;
			303: Pixel = 157;
			304: Pixel = 154;
			305: Pixel = 155;
			306: Pixel = 164;
			307: Pixel = 167;
			308: Pixel = 166;
			309: Pixel = 164;
			310: Pixel = 155;
			311: Pixel = 135;
			312: Pixel = 102;
			313: Pixel = 89;
			314: Pixel = 99;
			315: Pixel = 104;
			316: Pixel = 106;
			317: Pixel = 105;
			318: Pixel = 103;
			319: Pixel = 102;
			320: Pixel = 108;
			321: Pixel = 115;
			322: Pixel = 119;
			323: Pixel = 123;
			324: Pixel = 125;
			325: Pixel = 127;
			326: Pixel = 129;
			327: Pixel = 130;
			328: Pixel = 130;
			329: Pixel = 131;
			330: Pixel = 130;
			331: Pixel = 131;
			332: Pixel = 131;
			333: Pixel = 132;
			334: Pixel = 133;
			335: Pixel = 131;
			336: Pixel = 132;
			337: Pixel = 130;
			338: Pixel = 132;
			339: Pixel = 132;
			340: Pixel = 132;
			341: Pixel = 132;
			342: Pixel = 132;
			343: Pixel = 130;
			344: Pixel = 131;
			345: Pixel = 129;
			346: Pixel = 130;
			347: Pixel = 135;
			348: Pixel = 135;
			349: Pixel = 131;
			350: Pixel = 131;
			351: Pixel = 131;
			352: Pixel = 128;
			353: Pixel = 129;
			354: Pixel = 128;
			355: Pixel = 126;
			356: Pixel = 128;
			357: Pixel = 129;
			358: Pixel = 128;
			359: Pixel = 127;
			360: Pixel = 122;
			361: Pixel = 116;
			362: Pixel = 112;
			363: Pixel = 103;
			364: Pixel = 119;
			365: Pixel = 144;
			366: Pixel = 154;
			367: Pixel = 161;
			368: Pixel = 161;
			369: Pixel = 160;
			370: Pixel = 163;
			371: Pixel = 161;
			372: Pixel = 157;
			373: Pixel = 157;
			374: Pixel = 154;
			375: Pixel = 154;
			376: Pixel = 151;
			377: Pixel = 152;
			378: Pixel = 152;
			379: Pixel = 146;
			380: Pixel = 182;
			381: Pixel = 215;
			382: Pixel = 221;
			383: Pixel = 199;
			384: Pixel = 114;
			385: Pixel = 107;
			386: Pixel = 116;
			387: Pixel = 118;
			388: Pixel = 122;
			389: Pixel = 122;
			390: Pixel = 122;
			391: Pixel = 123;
			392: Pixel = 125;
			393: Pixel = 126;
			394: Pixel = 130;
			395: Pixel = 136;
			396: Pixel = 93;
			397: Pixel = 45;
			398: Pixel = 47;
			399: Pixel = 49;
			400: Pixel = 154;
			401: Pixel = 156;
			402: Pixel = 158;
			403: Pixel = 158;
			404: Pixel = 155;
			405: Pixel = 158;
			406: Pixel = 166;
			407: Pixel = 165;
			408: Pixel = 162;
			409: Pixel = 160;
			410: Pixel = 156;
			411: Pixel = 137;
			412: Pixel = 103;
			413: Pixel = 88;
			414: Pixel = 98;
			415: Pixel = 105;
			416: Pixel = 104;
			417: Pixel = 104;
			418: Pixel = 102;
			419: Pixel = 103;
			420: Pixel = 109;
			421: Pixel = 114;
			422: Pixel = 119;
			423: Pixel = 122;
			424: Pixel = 125;
			425: Pixel = 127;
			426: Pixel = 128;
			427: Pixel = 129;
			428: Pixel = 130;
			429: Pixel = 129;
			430: Pixel = 129;
			431: Pixel = 130;
			432: Pixel = 130;
			433: Pixel = 131;
			434: Pixel = 131;
			435: Pixel = 129;
			436: Pixel = 130;
			437: Pixel = 132;
			438: Pixel = 131;
			439: Pixel = 129;
			440: Pixel = 129;
			441: Pixel = 128;
			442: Pixel = 128;
			443: Pixel = 129;
			444: Pixel = 129;
			445: Pixel = 127;
			446: Pixel = 128;
			447: Pixel = 131;
			448: Pixel = 134;
			449: Pixel = 131;
			450: Pixel = 130;
			451: Pixel = 130;
			452: Pixel = 128;
			453: Pixel = 128;
			454: Pixel = 126;
			455: Pixel = 126;
			456: Pixel = 127;
			457: Pixel = 127;
			458: Pixel = 127;
			459: Pixel = 125;
			460: Pixel = 123;
			461: Pixel = 119;
			462: Pixel = 110;
			463: Pixel = 105;
			464: Pixel = 112;
			465: Pixel = 138;
			466: Pixel = 153;
			467: Pixel = 161;
			468: Pixel = 163;
			469: Pixel = 160;
			470: Pixel = 160;
			471: Pixel = 160;
			472: Pixel = 158;
			473: Pixel = 156;
			474: Pixel = 155;
			475: Pixel = 153;
			476: Pixel = 152;
			477: Pixel = 151;
			478: Pixel = 151;
			479: Pixel = 147;
			480: Pixel = 153;
			481: Pixel = 203;
			482: Pixel = 217;
			483: Pixel = 222;
			484: Pixel = 163;
			485: Pixel = 101;
			486: Pixel = 114;
			487: Pixel = 119;
			488: Pixel = 120;
			489: Pixel = 122;
			490: Pixel = 120;
			491: Pixel = 124;
			492: Pixel = 127;
			493: Pixel = 131;
			494: Pixel = 139;
			495: Pixel = 95;
			496: Pixel = 45;
			497: Pixel = 46;
			498: Pixel = 48;
			499: Pixel = 50;
			500: Pixel = 156;
			501: Pixel = 157;
			502: Pixel = 158;
			503: Pixel = 158;
			504: Pixel = 158;
			505: Pixel = 164;
			506: Pixel = 167;
			507: Pixel = 164;
			508: Pixel = 158;
			509: Pixel = 160;
			510: Pixel = 158;
			511: Pixel = 135;
			512: Pixel = 98;
			513: Pixel = 85;
			514: Pixel = 97;
			515: Pixel = 104;
			516: Pixel = 105;
			517: Pixel = 105;
			518: Pixel = 102;
			519: Pixel = 104;
			520: Pixel = 107;
			521: Pixel = 114;
			522: Pixel = 120;
			523: Pixel = 122;
			524: Pixel = 125;
			525: Pixel = 127;
			526: Pixel = 126;
			527: Pixel = 128;
			528: Pixel = 127;
			529: Pixel = 129;
			530: Pixel = 129;
			531: Pixel = 130;
			532: Pixel = 129;
			533: Pixel = 129;
			534: Pixel = 130;
			535: Pixel = 128;
			536: Pixel = 129;
			537: Pixel = 134;
			538: Pixel = 133;
			539: Pixel = 127;
			540: Pixel = 123;
			541: Pixel = 123;
			542: Pixel = 125;
			543: Pixel = 127;
			544: Pixel = 125;
			545: Pixel = 125;
			546: Pixel = 126;
			547: Pixel = 128;
			548: Pixel = 129;
			549: Pixel = 130;
			550: Pixel = 131;
			551: Pixel = 129;
			552: Pixel = 126;
			553: Pixel = 127;
			554: Pixel = 127;
			555: Pixel = 126;
			556: Pixel = 126;
			557: Pixel = 125;
			558: Pixel = 127;
			559: Pixel = 126;
			560: Pixel = 122;
			561: Pixel = 120;
			562: Pixel = 112;
			563: Pixel = 106;
			564: Pixel = 116;
			565: Pixel = 135;
			566: Pixel = 152;
			567: Pixel = 159;
			568: Pixel = 161;
			569: Pixel = 160;
			570: Pixel = 158;
			571: Pixel = 158;
			572: Pixel = 158;
			573: Pixel = 156;
			574: Pixel = 155;
			575: Pixel = 155;
			576: Pixel = 154;
			577: Pixel = 153;
			578: Pixel = 151;
			579: Pixel = 150;
			580: Pixel = 142;
			581: Pixel = 175;
			582: Pixel = 215;
			583: Pixel = 220;
			584: Pixel = 212;
			585: Pixel = 126;
			586: Pixel = 105;
			587: Pixel = 119;
			588: Pixel = 121;
			589: Pixel = 122;
			590: Pixel = 120;
			591: Pixel = 121;
			592: Pixel = 126;
			593: Pixel = 137;
			594: Pixel = 90;
			595: Pixel = 43;
			596: Pixel = 46;
			597: Pixel = 45;
			598: Pixel = 48;
			599: Pixel = 53;
			600: Pixel = 158;
			601: Pixel = 158;
			602: Pixel = 160;
			603: Pixel = 160;
			604: Pixel = 164;
			605: Pixel = 169;
			606: Pixel = 168;
			607: Pixel = 162;
			608: Pixel = 157;
			609: Pixel = 160;
			610: Pixel = 159;
			611: Pixel = 135;
			612: Pixel = 100;
			613: Pixel = 89;
			614: Pixel = 98;
			615: Pixel = 103;
			616: Pixel = 106;
			617: Pixel = 104;
			618: Pixel = 102;
			619: Pixel = 103;
			620: Pixel = 107;
			621: Pixel = 114;
			622: Pixel = 119;
			623: Pixel = 122;
			624: Pixel = 123;
			625: Pixel = 126;
			626: Pixel = 127;
			627: Pixel = 128;
			628: Pixel = 127;
			629: Pixel = 127;
			630: Pixel = 129;
			631: Pixel = 130;
			632: Pixel = 129;
			633: Pixel = 129;
			634: Pixel = 129;
			635: Pixel = 130;
			636: Pixel = 128;
			637: Pixel = 131;
			638: Pixel = 131;
			639: Pixel = 126;
			640: Pixel = 123;
			641: Pixel = 122;
			642: Pixel = 122;
			643: Pixel = 126;
			644: Pixel = 126;
			645: Pixel = 124;
			646: Pixel = 124;
			647: Pixel = 128;
			648: Pixel = 129;
			649: Pixel = 129;
			650: Pixel = 132;
			651: Pixel = 128;
			652: Pixel = 127;
			653: Pixel = 128;
			654: Pixel = 127;
			655: Pixel = 126;
			656: Pixel = 126;
			657: Pixel = 126;
			658: Pixel = 127;
			659: Pixel = 127;
			660: Pixel = 123;
			661: Pixel = 118;
			662: Pixel = 112;
			663: Pixel = 107;
			664: Pixel = 115;
			665: Pixel = 133;
			666: Pixel = 147;
			667: Pixel = 155;
			668: Pixel = 159;
			669: Pixel = 158;
			670: Pixel = 157;
			671: Pixel = 159;
			672: Pixel = 157;
			673: Pixel = 156;
			674: Pixel = 156;
			675: Pixel = 156;
			676: Pixel = 155;
			677: Pixel = 155;
			678: Pixel = 153;
			679: Pixel = 152;
			680: Pixel = 146;
			681: Pixel = 146;
			682: Pixel = 196;
			683: Pixel = 217;
			684: Pixel = 225;
			685: Pixel = 187;
			686: Pixel = 107;
			687: Pixel = 111;
			688: Pixel = 118;
			689: Pixel = 122;
			690: Pixel = 122;
			691: Pixel = 126;
			692: Pixel = 135;
			693: Pixel = 92;
			694: Pixel = 40;
			695: Pixel = 47;
			696: Pixel = 50;
			697: Pixel = 51;
			698: Pixel = 50;
			699: Pixel = 53;
			700: Pixel = 159;
			701: Pixel = 160;
			702: Pixel = 161;
			703: Pixel = 164;
			704: Pixel = 168;
			705: Pixel = 165;
			706: Pixel = 164;
			707: Pixel = 160;
			708: Pixel = 158;
			709: Pixel = 161;
			710: Pixel = 156;
			711: Pixel = 134;
			712: Pixel = 96;
			713: Pixel = 84;
			714: Pixel = 97;
			715: Pixel = 103;
			716: Pixel = 102;
			717: Pixel = 102;
			718: Pixel = 102;
			719: Pixel = 102;
			720: Pixel = 107;
			721: Pixel = 114;
			722: Pixel = 118;
			723: Pixel = 119;
			724: Pixel = 122;
			725: Pixel = 124;
			726: Pixel = 125;
			727: Pixel = 127;
			728: Pixel = 125;
			729: Pixel = 124;
			730: Pixel = 127;
			731: Pixel = 129;
			732: Pixel = 127;
			733: Pixel = 127;
			734: Pixel = 129;
			735: Pixel = 130;
			736: Pixel = 128;
			737: Pixel = 129;
			738: Pixel = 128;
			739: Pixel = 126;
			740: Pixel = 125;
			741: Pixel = 123;
			742: Pixel = 123;
			743: Pixel = 121;
			744: Pixel = 119;
			745: Pixel = 117;
			746: Pixel = 120;
			747: Pixel = 125;
			748: Pixel = 129;
			749: Pixel = 130;
			750: Pixel = 131;
			751: Pixel = 127;
			752: Pixel = 126;
			753: Pixel = 128;
			754: Pixel = 127;
			755: Pixel = 125;
			756: Pixel = 125;
			757: Pixel = 126;
			758: Pixel = 126;
			759: Pixel = 126;
			760: Pixel = 121;
			761: Pixel = 118;
			762: Pixel = 116;
			763: Pixel = 109;
			764: Pixel = 114;
			765: Pixel = 131;
			766: Pixel = 144;
			767: Pixel = 151;
			768: Pixel = 155;
			769: Pixel = 157;
			770: Pixel = 156;
			771: Pixel = 157;
			772: Pixel = 155;
			773: Pixel = 156;
			774: Pixel = 154;
			775: Pixel = 156;
			776: Pixel = 156;
			777: Pixel = 154;
			778: Pixel = 153;
			779: Pixel = 150;
			780: Pixel = 148;
			781: Pixel = 138;
			782: Pixel = 166;
			783: Pixel = 216;
			784: Pixel = 221;
			785: Pixel = 222;
			786: Pixel = 144;
			787: Pixel = 99;
			788: Pixel = 114;
			789: Pixel = 118;
			790: Pixel = 124;
			791: Pixel = 135;
			792: Pixel = 90;
			793: Pixel = 40;
			794: Pixel = 43;
			795: Pixel = 53;
			796: Pixel = 56;
			797: Pixel = 52;
			798: Pixel = 49;
			799: Pixel = 47;
			800: Pixel = 161;
			801: Pixel = 160;
			802: Pixel = 162;
			803: Pixel = 168;
			804: Pixel = 162;
			805: Pixel = 157;
			806: Pixel = 157;
			807: Pixel = 160;
			808: Pixel = 159;
			809: Pixel = 161;
			810: Pixel = 157;
			811: Pixel = 134;
			812: Pixel = 95;
			813: Pixel = 84;
			814: Pixel = 97;
			815: Pixel = 103;
			816: Pixel = 103;
			817: Pixel = 103;
			818: Pixel = 102;
			819: Pixel = 102;
			820: Pixel = 106;
			821: Pixel = 114;
			822: Pixel = 119;
			823: Pixel = 120;
			824: Pixel = 123;
			825: Pixel = 123;
			826: Pixel = 125;
			827: Pixel = 125;
			828: Pixel = 124;
			829: Pixel = 126;
			830: Pixel = 128;
			831: Pixel = 127;
			832: Pixel = 126;
			833: Pixel = 129;
			834: Pixel = 129;
			835: Pixel = 128;
			836: Pixel = 128;
			837: Pixel = 129;
			838: Pixel = 126;
			839: Pixel = 124;
			840: Pixel = 127;
			841: Pixel = 124;
			842: Pixel = 123;
			843: Pixel = 130;
			844: Pixel = 131;
			845: Pixel = 127;
			846: Pixel = 122;
			847: Pixel = 117;
			848: Pixel = 119;
			849: Pixel = 124;
			850: Pixel = 128;
			851: Pixel = 127;
			852: Pixel = 126;
			853: Pixel = 127;
			854: Pixel = 129;
			855: Pixel = 127;
			856: Pixel = 127;
			857: Pixel = 126;
			858: Pixel = 126;
			859: Pixel = 125;
			860: Pixel = 121;
			861: Pixel = 116;
			862: Pixel = 115;
			863: Pixel = 109;
			864: Pixel = 113;
			865: Pixel = 129;
			866: Pixel = 142;
			867: Pixel = 147;
			868: Pixel = 151;
			869: Pixel = 155;
			870: Pixel = 156;
			871: Pixel = 154;
			872: Pixel = 154;
			873: Pixel = 154;
			874: Pixel = 153;
			875: Pixel = 154;
			876: Pixel = 155;
			877: Pixel = 152;
			878: Pixel = 148;
			879: Pixel = 146;
			880: Pixel = 144;
			881: Pixel = 141;
			882: Pixel = 142;
			883: Pixel = 194;
			884: Pixel = 220;
			885: Pixel = 226;
			886: Pixel = 198;
			887: Pixel = 109;
			888: Pixel = 106;
			889: Pixel = 114;
			890: Pixel = 128;
			891: Pixel = 93;
			892: Pixel = 42;
			893: Pixel = 44;
			894: Pixel = 50;
			895: Pixel = 57;
			896: Pixel = 55;
			897: Pixel = 51;
			898: Pixel = 46;
			899: Pixel = 45;
			900: Pixel = 162;
			901: Pixel = 159;
			902: Pixel = 167;
			903: Pixel = 166;
			904: Pixel = 152;
			905: Pixel = 147;
			906: Pixel = 151;
			907: Pixel = 162;
			908: Pixel = 160;
			909: Pixel = 162;
			910: Pixel = 158;
			911: Pixel = 136;
			912: Pixel = 98;
			913: Pixel = 85;
			914: Pixel = 96;
			915: Pixel = 102;
			916: Pixel = 105;
			917: Pixel = 103;
			918: Pixel = 103;
			919: Pixel = 103;
			920: Pixel = 110;
			921: Pixel = 113;
			922: Pixel = 119;
			923: Pixel = 121;
			924: Pixel = 123;
			925: Pixel = 124;
			926: Pixel = 125;
			927: Pixel = 126;
			928: Pixel = 126;
			929: Pixel = 129;
			930: Pixel = 129;
			931: Pixel = 128;
			932: Pixel = 127;
			933: Pixel = 129;
			934: Pixel = 130;
			935: Pixel = 128;
			936: Pixel = 125;
			937: Pixel = 127;
			938: Pixel = 135;
			939: Pixel = 137;
			940: Pixel = 142;
			941: Pixel = 147;
			942: Pixel = 157;
			943: Pixel = 172;
			944: Pixel = 176;
			945: Pixel = 177;
			946: Pixel = 176;
			947: Pixel = 164;
			948: Pixel = 147;
			949: Pixel = 125;
			950: Pixel = 114;
			951: Pixel = 120;
			952: Pixel = 125;
			953: Pixel = 129;
			954: Pixel = 130;
			955: Pixel = 128;
			956: Pixel = 126;
			957: Pixel = 126;
			958: Pixel = 126;
			959: Pixel = 125;
			960: Pixel = 121;
			961: Pixel = 117;
			962: Pixel = 113;
			963: Pixel = 108;
			964: Pixel = 111;
			965: Pixel = 128;
			966: Pixel = 141;
			967: Pixel = 144;
			968: Pixel = 146;
			969: Pixel = 151;
			970: Pixel = 154;
			971: Pixel = 154;
			972: Pixel = 152;
			973: Pixel = 153;
			974: Pixel = 154;
			975: Pixel = 153;
			976: Pixel = 151;
			977: Pixel = 149;
			978: Pixel = 145;
			979: Pixel = 144;
			980: Pixel = 142;
			981: Pixel = 143;
			982: Pixel = 138;
			983: Pixel = 161;
			984: Pixel = 212;
			985: Pixel = 221;
			986: Pixel = 225;
			987: Pixel = 159;
			988: Pixel = 103;
			989: Pixel = 124;
			990: Pixel = 88;
			991: Pixel = 40;
			992: Pixel = 43;
			993: Pixel = 47;
			994: Pixel = 53;
			995: Pixel = 58;
			996: Pixel = 55;
			997: Pixel = 45;
			998: Pixel = 45;
			999: Pixel = 47;
			1000: Pixel = 159;
			1001: Pixel = 162;
			1002: Pixel = 169;
			1003: Pixel = 160;
			1004: Pixel = 141;
			1005: Pixel = 134;
			1006: Pixel = 149;
			1007: Pixel = 164;
			1008: Pixel = 161;
			1009: Pixel = 164;
			1010: Pixel = 158;
			1011: Pixel = 136;
			1012: Pixel = 96;
			1013: Pixel = 83;
			1014: Pixel = 94;
			1015: Pixel = 100;
			1016: Pixel = 102;
			1017: Pixel = 102;
			1018: Pixel = 104;
			1019: Pixel = 104;
			1020: Pixel = 110;
			1021: Pixel = 116;
			1022: Pixel = 120;
			1023: Pixel = 121;
			1024: Pixel = 124;
			1025: Pixel = 126;
			1026: Pixel = 124;
			1027: Pixel = 126;
			1028: Pixel = 129;
			1029: Pixel = 128;
			1030: Pixel = 129;
			1031: Pixel = 127;
			1032: Pixel = 123;
			1033: Pixel = 125;
			1034: Pixel = 129;
			1035: Pixel = 127;
			1036: Pixel = 131;
			1037: Pixel = 141;
			1038: Pixel = 150;
			1039: Pixel = 146;
			1040: Pixel = 147;
			1041: Pixel = 160;
			1042: Pixel = 166;
			1043: Pixel = 170;
			1044: Pixel = 181;
			1045: Pixel = 176;
			1046: Pixel = 174;
			1047: Pixel = 184;
			1048: Pixel = 190;
			1049: Pixel = 187;
			1050: Pixel = 166;
			1051: Pixel = 128;
			1052: Pixel = 112;
			1053: Pixel = 123;
			1054: Pixel = 128;
			1055: Pixel = 127;
			1056: Pixel = 126;
			1057: Pixel = 125;
			1058: Pixel = 124;
			1059: Pixel = 122;
			1060: Pixel = 118;
			1061: Pixel = 115;
			1062: Pixel = 113;
			1063: Pixel = 108;
			1064: Pixel = 111;
			1065: Pixel = 130;
			1066: Pixel = 143;
			1067: Pixel = 144;
			1068: Pixel = 144;
			1069: Pixel = 148;
			1070: Pixel = 152;
			1071: Pixel = 153;
			1072: Pixel = 151;
			1073: Pixel = 151;
			1074: Pixel = 149;
			1075: Pixel = 149;
			1076: Pixel = 147;
			1077: Pixel = 144;
			1078: Pixel = 143;
			1079: Pixel = 140;
			1080: Pixel = 140;
			1081: Pixel = 141;
			1082: Pixel = 141;
			1083: Pixel = 138;
			1084: Pixel = 183;
			1085: Pixel = 220;
			1086: Pixel = 226;
			1087: Pixel = 213;
			1088: Pixel = 137;
			1089: Pixel = 90;
			1090: Pixel = 41;
			1091: Pixel = 43;
			1092: Pixel = 48;
			1093: Pixel = 51;
			1094: Pixel = 53;
			1095: Pixel = 51;
			1096: Pixel = 48;
			1097: Pixel = 48;
			1098: Pixel = 46;
			1099: Pixel = 45;
			1100: Pixel = 160;
			1101: Pixel = 169;
			1102: Pixel = 166;
			1103: Pixel = 148;
			1104: Pixel = 122;
			1105: Pixel = 125;
			1106: Pixel = 154;
			1107: Pixel = 165;
			1108: Pixel = 164;
			1109: Pixel = 164;
			1110: Pixel = 159;
			1111: Pixel = 137;
			1112: Pixel = 94;
			1113: Pixel = 80;
			1114: Pixel = 93;
			1115: Pixel = 97;
			1116: Pixel = 100;
			1117: Pixel = 100;
			1118: Pixel = 100;
			1119: Pixel = 104;
			1120: Pixel = 108;
			1121: Pixel = 115;
			1122: Pixel = 118;
			1123: Pixel = 121;
			1124: Pixel = 122;
			1125: Pixel = 123;
			1126: Pixel = 123;
			1127: Pixel = 125;
			1128: Pixel = 126;
			1129: Pixel = 127;
			1130: Pixel = 124;
			1131: Pixel = 126;
			1132: Pixel = 136;
			1133: Pixel = 142;
			1134: Pixel = 137;
			1135: Pixel = 123;
			1136: Pixel = 133;
			1137: Pixel = 140;
			1138: Pixel = 138;
			1139: Pixel = 144;
			1140: Pixel = 148;
			1141: Pixel = 151;
			1142: Pixel = 158;
			1143: Pixel = 165;
			1144: Pixel = 169;
			1145: Pixel = 174;
			1146: Pixel = 176;
			1147: Pixel = 179;
			1148: Pixel = 184;
			1149: Pixel = 190;
			1150: Pixel = 200;
			1151: Pixel = 194;
			1152: Pixel = 151;
			1153: Pixel = 113;
			1154: Pixel = 118;
			1155: Pixel = 126;
			1156: Pixel = 122;
			1157: Pixel = 123;
			1158: Pixel = 122;
			1159: Pixel = 119;
			1160: Pixel = 115;
			1161: Pixel = 113;
			1162: Pixel = 110;
			1163: Pixel = 105;
			1164: Pixel = 111;
			1165: Pixel = 129;
			1166: Pixel = 143;
			1167: Pixel = 146;
			1168: Pixel = 144;
			1169: Pixel = 147;
			1170: Pixel = 148;
			1171: Pixel = 151;
			1172: Pixel = 151;
			1173: Pixel = 147;
			1174: Pixel = 145;
			1175: Pixel = 145;
			1176: Pixel = 146;
			1177: Pixel = 143;
			1178: Pixel = 142;
			1179: Pixel = 140;
			1180: Pixel = 139;
			1181: Pixel = 140;
			1182: Pixel = 142;
			1183: Pixel = 137;
			1184: Pixel = 146;
			1185: Pixel = 207;
			1186: Pixel = 221;
			1187: Pixel = 236;
			1188: Pixel = 174;
			1189: Pixel = 38;
			1190: Pixel = 42;
			1191: Pixel = 46;
			1192: Pixel = 52;
			1193: Pixel = 54;
			1194: Pixel = 53;
			1195: Pixel = 48;
			1196: Pixel = 51;
			1197: Pixel = 51;
			1198: Pixel = 46;
			1199: Pixel = 48;
			1200: Pixel = 168;
			1201: Pixel = 171;
			1202: Pixel = 158;
			1203: Pixel = 132;
			1204: Pixel = 94;
			1205: Pixel = 123;
			1206: Pixel = 157;
			1207: Pixel = 166;
			1208: Pixel = 165;
			1209: Pixel = 164;
			1210: Pixel = 159;
			1211: Pixel = 137;
			1212: Pixel = 94;
			1213: Pixel = 77;
			1214: Pixel = 87;
			1215: Pixel = 95;
			1216: Pixel = 96;
			1217: Pixel = 98;
			1218: Pixel = 100;
			1219: Pixel = 103;
			1220: Pixel = 106;
			1221: Pixel = 111;
			1222: Pixel = 116;
			1223: Pixel = 118;
			1224: Pixel = 119;
			1225: Pixel = 123;
			1226: Pixel = 122;
			1227: Pixel = 124;
			1228: Pixel = 125;
			1229: Pixel = 122;
			1230: Pixel = 134;
			1231: Pixel = 130;
			1232: Pixel = 131;
			1233: Pixel = 129;
			1234: Pixel = 122;
			1235: Pixel = 121;
			1236: Pixel = 129;
			1237: Pixel = 131;
			1238: Pixel = 129;
			1239: Pixel = 137;
			1240: Pixel = 143;
			1241: Pixel = 149;
			1242: Pixel = 157;
			1243: Pixel = 160;
			1244: Pixel = 168;
			1245: Pixel = 174;
			1246: Pixel = 183;
			1247: Pixel = 185;
			1248: Pixel = 185;
			1249: Pixel = 187;
			1250: Pixel = 188;
			1251: Pixel = 196;
			1252: Pixel = 202;
			1253: Pixel = 176;
			1254: Pixel = 122;
			1255: Pixel = 105;
			1256: Pixel = 119;
			1257: Pixel = 120;
			1258: Pixel = 119;
			1259: Pixel = 118;
			1260: Pixel = 115;
			1261: Pixel = 111;
			1262: Pixel = 108;
			1263: Pixel = 102;
			1264: Pixel = 108;
			1265: Pixel = 129;
			1266: Pixel = 144;
			1267: Pixel = 148;
			1268: Pixel = 144;
			1269: Pixel = 145;
			1270: Pixel = 146;
			1271: Pixel = 146;
			1272: Pixel = 150;
			1273: Pixel = 148;
			1274: Pixel = 141;
			1275: Pixel = 141;
			1276: Pixel = 144;
			1277: Pixel = 144;
			1278: Pixel = 143;
			1279: Pixel = 142;
			1280: Pixel = 140;
			1281: Pixel = 140;
			1282: Pixel = 143;
			1283: Pixel = 143;
			1284: Pixel = 137;
			1285: Pixel = 169;
			1286: Pixel = 223;
			1287: Pixel = 236;
			1288: Pixel = 110;
			1289: Pixel = 30;
			1290: Pixel = 46;
			1291: Pixel = 50;
			1292: Pixel = 54;
			1293: Pixel = 54;
			1294: Pixel = 45;
			1295: Pixel = 46;
			1296: Pixel = 52;
			1297: Pixel = 43;
			1298: Pixel = 49;
			1299: Pixel = 52;
			1300: Pixel = 172;
			1301: Pixel = 165;
			1302: Pixel = 148;
			1303: Pixel = 104;
			1304: Pixel = 79;
			1305: Pixel = 124;
			1306: Pixel = 155;
			1307: Pixel = 167;
			1308: Pixel = 164;
			1309: Pixel = 164;
			1310: Pixel = 156;
			1311: Pixel = 134;
			1312: Pixel = 92;
			1313: Pixel = 74;
			1314: Pixel = 88;
			1315: Pixel = 95;
			1316: Pixel = 99;
			1317: Pixel = 99;
			1318: Pixel = 100;
			1319: Pixel = 101;
			1320: Pixel = 104;
			1321: Pixel = 110;
			1322: Pixel = 114;
			1323: Pixel = 114;
			1324: Pixel = 117;
			1325: Pixel = 120;
			1326: Pixel = 121;
			1327: Pixel = 124;
			1328: Pixel = 124;
			1329: Pixel = 121;
			1330: Pixel = 133;
			1331: Pixel = 112;
			1332: Pixel = 116;
			1333: Pixel = 118;
			1334: Pixel = 122;
			1335: Pixel = 121;
			1336: Pixel = 130;
			1337: Pixel = 130;
			1338: Pixel = 131;
			1339: Pixel = 135;
			1340: Pixel = 134;
			1341: Pixel = 140;
			1342: Pixel = 149;
			1343: Pixel = 161;
			1344: Pixel = 174;
			1345: Pixel = 175;
			1346: Pixel = 180;
			1347: Pixel = 182;
			1348: Pixel = 186;
			1349: Pixel = 189;
			1350: Pixel = 190;
			1351: Pixel = 194;
			1352: Pixel = 195;
			1353: Pixel = 199;
			1354: Pixel = 198;
			1355: Pixel = 141;
			1356: Pixel = 96;
			1357: Pixel = 103;
			1358: Pixel = 113;
			1359: Pixel = 114;
			1360: Pixel = 113;
			1361: Pixel = 109;
			1362: Pixel = 108;
			1363: Pixel = 103;
			1364: Pixel = 107;
			1365: Pixel = 129;
			1366: Pixel = 147;
			1367: Pixel = 151;
			1368: Pixel = 148;
			1369: Pixel = 144;
			1370: Pixel = 141;
			1371: Pixel = 140;
			1372: Pixel = 142;
			1373: Pixel = 149;
			1374: Pixel = 143;
			1375: Pixel = 141;
			1376: Pixel = 144;
			1377: Pixel = 144;
			1378: Pixel = 142;
			1379: Pixel = 142;
			1380: Pixel = 142;
			1381: Pixel = 143;
			1382: Pixel = 143;
			1383: Pixel = 144;
			1384: Pixel = 145;
			1385: Pixel = 148;
			1386: Pixel = 206;
			1387: Pixel = 133;
			1388: Pixel = 35;
			1389: Pixel = 44;
			1390: Pixel = 46;
			1391: Pixel = 51;
			1392: Pixel = 54;
			1393: Pixel = 50;
			1394: Pixel = 48;
			1395: Pixel = 52;
			1396: Pixel = 45;
			1397: Pixel = 52;
			1398: Pixel = 57;
			1399: Pixel = 29;
			1400: Pixel = 170;
			1401: Pixel = 158;
			1402: Pixel = 127;
			1403: Pixel = 81;
			1404: Pixel = 84;
			1405: Pixel = 125;
			1406: Pixel = 154;
			1407: Pixel = 168;
			1408: Pixel = 166;
			1409: Pixel = 163;
			1410: Pixel = 156;
			1411: Pixel = 135;
			1412: Pixel = 90;
			1413: Pixel = 74;
			1414: Pixel = 89;
			1415: Pixel = 97;
			1416: Pixel = 100;
			1417: Pixel = 100;
			1418: Pixel = 99;
			1419: Pixel = 100;
			1420: Pixel = 105;
			1421: Pixel = 110;
			1422: Pixel = 113;
			1423: Pixel = 114;
			1424: Pixel = 117;
			1425: Pixel = 119;
			1426: Pixel = 120;
			1427: Pixel = 123;
			1428: Pixel = 120;
			1429: Pixel = 137;
			1430: Pixel = 122;
			1431: Pixel = 111;
			1432: Pixel = 112;
			1433: Pixel = 116;
			1434: Pixel = 122;
			1435: Pixel = 126;
			1436: Pixel = 127;
			1437: Pixel = 131;
			1438: Pixel = 136;
			1439: Pixel = 135;
			1440: Pixel = 136;
			1441: Pixel = 138;
			1442: Pixel = 146;
			1443: Pixel = 155;
			1444: Pixel = 164;
			1445: Pixel = 172;
			1446: Pixel = 180;
			1447: Pixel = 183;
			1448: Pixel = 189;
			1449: Pixel = 191;
			1450: Pixel = 193;
			1451: Pixel = 197;
			1452: Pixel = 195;
			1453: Pixel = 192;
			1454: Pixel = 196;
			1455: Pixel = 204;
			1456: Pixel = 159;
			1457: Pixel = 112;
			1458: Pixel = 95;
			1459: Pixel = 111;
			1460: Pixel = 109;
			1461: Pixel = 105;
			1462: Pixel = 107;
			1463: Pixel = 102;
			1464: Pixel = 105;
			1465: Pixel = 130;
			1466: Pixel = 150;
			1467: Pixel = 155;
			1468: Pixel = 153;
			1469: Pixel = 148;
			1470: Pixel = 135;
			1471: Pixel = 127;
			1472: Pixel = 129;
			1473: Pixel = 145;
			1474: Pixel = 147;
			1475: Pixel = 142;
			1476: Pixel = 146;
			1477: Pixel = 145;
			1478: Pixel = 142;
			1479: Pixel = 142;
			1480: Pixel = 144;
			1481: Pixel = 144;
			1482: Pixel = 145;
			1483: Pixel = 147;
			1484: Pixel = 148;
			1485: Pixel = 161;
			1486: Pixel = 110;
			1487: Pixel = 37;
			1488: Pixel = 43;
			1489: Pixel = 46;
			1490: Pixel = 53;
			1491: Pixel = 52;
			1492: Pixel = 46;
			1493: Pixel = 46;
			1494: Pixel = 56;
			1495: Pixel = 48;
			1496: Pixel = 51;
			1497: Pixel = 65;
			1498: Pixel = 37;
			1499: Pixel = 75;
			1500: Pixel = 162;
			1501: Pixel = 145;
			1502: Pixel = 99;
			1503: Pixel = 79;
			1504: Pixel = 88;
			1505: Pixel = 126;
			1506: Pixel = 154;
			1507: Pixel = 166;
			1508: Pixel = 167;
			1509: Pixel = 164;
			1510: Pixel = 157;
			1511: Pixel = 134;
			1512: Pixel = 90;
			1513: Pixel = 75;
			1514: Pixel = 89;
			1515: Pixel = 98;
			1516: Pixel = 99;
			1517: Pixel = 99;
			1518: Pixel = 100;
			1519: Pixel = 101;
			1520: Pixel = 105;
			1521: Pixel = 110;
			1522: Pixel = 114;
			1523: Pixel = 114;
			1524: Pixel = 118;
			1525: Pixel = 121;
			1526: Pixel = 121;
			1527: Pixel = 120;
			1528: Pixel = 124;
			1529: Pixel = 133;
			1530: Pixel = 112;
			1531: Pixel = 107;
			1532: Pixel = 114;
			1533: Pixel = 117;
			1534: Pixel = 119;
			1535: Pixel = 124;
			1536: Pixel = 125;
			1537: Pixel = 127;
			1538: Pixel = 129;
			1539: Pixel = 135;
			1540: Pixel = 134;
			1541: Pixel = 137;
			1542: Pixel = 145;
			1543: Pixel = 150;
			1544: Pixel = 162;
			1545: Pixel = 178;
			1546: Pixel = 185;
			1547: Pixel = 184;
			1548: Pixel = 186;
			1549: Pixel = 192;
			1550: Pixel = 191;
			1551: Pixel = 188;
			1552: Pixel = 189;
			1553: Pixel = 196;
			1554: Pixel = 204;
			1555: Pixel = 211;
			1556: Pixel = 227;
			1557: Pixel = 224;
			1558: Pixel = 110;
			1559: Pixel = 90;
			1560: Pixel = 107;
			1561: Pixel = 101;
			1562: Pixel = 103;
			1563: Pixel = 99;
			1564: Pixel = 105;
			1565: Pixel = 130;
			1566: Pixel = 150;
			1567: Pixel = 155;
			1568: Pixel = 154;
			1569: Pixel = 152;
			1570: Pixel = 135;
			1571: Pixel = 107;
			1572: Pixel = 107;
			1573: Pixel = 133;
			1574: Pixel = 148;
			1575: Pixel = 145;
			1576: Pixel = 145;
			1577: Pixel = 145;
			1578: Pixel = 142;
			1579: Pixel = 143;
			1580: Pixel = 144;
			1581: Pixel = 144;
			1582: Pixel = 146;
			1583: Pixel = 146;
			1584: Pixel = 157;
			1585: Pixel = 130;
			1586: Pixel = 46;
			1587: Pixel = 43;
			1588: Pixel = 45;
			1589: Pixel = 49;
			1590: Pixel = 53;
			1591: Pixel = 48;
			1592: Pixel = 45;
			1593: Pixel = 55;
			1594: Pixel = 48;
			1595: Pixel = 46;
			1596: Pixel = 70;
			1597: Pixel = 52;
			1598: Pixel = 64;
			1599: Pixel = 155;
			1600: Pixel = 153;
			1601: Pixel = 119;
			1602: Pixel = 83;
			1603: Pixel = 84;
			1604: Pixel = 90;
			1605: Pixel = 125;
			1606: Pixel = 154;
			1607: Pixel = 166;
			1608: Pixel = 167;
			1609: Pixel = 165;
			1610: Pixel = 155;
			1611: Pixel = 131;
			1612: Pixel = 92;
			1613: Pixel = 76;
			1614: Pixel = 90;
			1615: Pixel = 96;
			1616: Pixel = 99;
			1617: Pixel = 100;
			1618: Pixel = 102;
			1619: Pixel = 101;
			1620: Pixel = 104;
			1621: Pixel = 111;
			1622: Pixel = 113;
			1623: Pixel = 115;
			1624: Pixel = 118;
			1625: Pixel = 121;
			1626: Pixel = 121;
			1627: Pixel = 122;
			1628: Pixel = 127;
			1629: Pixel = 111;
			1630: Pixel = 107;
			1631: Pixel = 114;
			1632: Pixel = 119;
			1633: Pixel = 119;
			1634: Pixel = 121;
			1635: Pixel = 119;
			1636: Pixel = 120;
			1637: Pixel = 127;
			1638: Pixel = 133;
			1639: Pixel = 135;
			1640: Pixel = 133;
			1641: Pixel = 137;
			1642: Pixel = 139;
			1643: Pixel = 151;
			1644: Pixel = 162;
			1645: Pixel = 177;
			1646: Pixel = 183;
			1647: Pixel = 189;
			1648: Pixel = 186;
			1649: Pixel = 178;
			1650: Pixel = 184;
			1651: Pixel = 197;
			1652: Pixel = 207;
			1653: Pixel = 211;
			1654: Pixel = 210;
			1655: Pixel = 210;
			1656: Pixel = 207;
			1657: Pixel = 228;
			1658: Pixel = 195;
			1659: Pixel = 83;
			1660: Pixel = 93;
			1661: Pixel = 100;
			1662: Pixel = 99;
			1663: Pixel = 96;
			1664: Pixel = 102;
			1665: Pixel = 128;
			1666: Pixel = 148;
			1667: Pixel = 154;
			1668: Pixel = 152;
			1669: Pixel = 152;
			1670: Pixel = 140;
			1671: Pixel = 97;
			1672: Pixel = 69;
			1673: Pixel = 111;
			1674: Pixel = 142;
			1675: Pixel = 147;
			1676: Pixel = 144;
			1677: Pixel = 145;
			1678: Pixel = 143;
			1679: Pixel = 143;
			1680: Pixel = 144;
			1681: Pixel = 144;
			1682: Pixel = 144;
			1683: Pixel = 152;
			1684: Pixel = 149;
			1685: Pixel = 60;
			1686: Pixel = 36;
			1687: Pixel = 44;
			1688: Pixel = 51;
			1689: Pixel = 54;
			1690: Pixel = 50;
			1691: Pixel = 44;
			1692: Pixel = 53;
			1693: Pixel = 49;
			1694: Pixel = 48;
			1695: Pixel = 62;
			1696: Pixel = 69;
			1697: Pixel = 72;
			1698: Pixel = 138;
			1699: Pixel = 156;
			1700: Pixel = 134;
			1701: Pixel = 92;
			1702: Pixel = 85;
			1703: Pixel = 88;
			1704: Pixel = 89;
			1705: Pixel = 125;
			1706: Pixel = 153;
			1707: Pixel = 166;
			1708: Pixel = 166;
			1709: Pixel = 165;
			1710: Pixel = 155;
			1711: Pixel = 131;
			1712: Pixel = 92;
			1713: Pixel = 77;
			1714: Pixel = 90;
			1715: Pixel = 95;
			1716: Pixel = 98;
			1717: Pixel = 102;
			1718: Pixel = 102;
			1719: Pixel = 100;
			1720: Pixel = 105;
			1721: Pixel = 109;
			1722: Pixel = 114;
			1723: Pixel = 116;
			1724: Pixel = 119;
			1725: Pixel = 121;
			1726: Pixel = 121;
			1727: Pixel = 125;
			1728: Pixel = 114;
			1729: Pixel = 106;
			1730: Pixel = 111;
			1731: Pixel = 115;
			1732: Pixel = 119;
			1733: Pixel = 118;
			1734: Pixel = 115;
			1735: Pixel = 117;
			1736: Pixel = 124;
			1737: Pixel = 129;
			1738: Pixel = 137;
			1739: Pixel = 136;
			1740: Pixel = 138;
			1741: Pixel = 142;
			1742: Pixel = 144;
			1743: Pixel = 148;
			1744: Pixel = 158;
			1745: Pixel = 174;
			1746: Pixel = 181;
			1747: Pixel = 173;
			1748: Pixel = 172;
			1749: Pixel = 190;
			1750: Pixel = 209;
			1751: Pixel = 210;
			1752: Pixel = 205;
			1753: Pixel = 205;
			1754: Pixel = 205;
			1755: Pixel = 205;
			1756: Pixel = 208;
			1757: Pixel = 211;
			1758: Pixel = 232;
			1759: Pixel = 166;
			1760: Pixel = 71;
			1761: Pixel = 91;
			1762: Pixel = 97;
			1763: Pixel = 94;
			1764: Pixel = 101;
			1765: Pixel = 127;
			1766: Pixel = 149;
			1767: Pixel = 155;
			1768: Pixel = 153;
			1769: Pixel = 151;
			1770: Pixel = 143;
			1771: Pixel = 104;
			1772: Pixel = 47;
			1773: Pixel = 80;
			1774: Pixel = 127;
			1775: Pixel = 147;
			1776: Pixel = 146;
			1777: Pixel = 144;
			1778: Pixel = 143;
			1779: Pixel = 143;
			1780: Pixel = 144;
			1781: Pixel = 143;
			1782: Pixel = 146;
			1783: Pixel = 157;
			1784: Pixel = 90;
			1785: Pixel = 43;
			1786: Pixel = 45;
			1787: Pixel = 50;
			1788: Pixel = 55;
			1789: Pixel = 54;
			1790: Pixel = 45;
			1791: Pixel = 53;
			1792: Pixel = 51;
			1793: Pixel = 45;
			1794: Pixel = 60;
			1795: Pixel = 71;
			1796: Pixel = 80;
			1797: Pixel = 133;
			1798: Pixel = 152;
			1799: Pixel = 139;
			1800: Pixel = 103;
			1801: Pixel = 84;
			1802: Pixel = 92;
			1803: Pixel = 88;
			1804: Pixel = 88;
			1805: Pixel = 123;
			1806: Pixel = 151;
			1807: Pixel = 164;
			1808: Pixel = 167;
			1809: Pixel = 164;
			1810: Pixel = 156;
			1811: Pixel = 131;
			1812: Pixel = 91;
			1813: Pixel = 77;
			1814: Pixel = 93;
			1815: Pixel = 99;
			1816: Pixel = 98;
			1817: Pixel = 99;
			1818: Pixel = 100;
			1819: Pixel = 101;
			1820: Pixel = 104;
			1821: Pixel = 109;
			1822: Pixel = 115;
			1823: Pixel = 117;
			1824: Pixel = 118;
			1825: Pixel = 120;
			1826: Pixel = 124;
			1827: Pixel = 120;
			1828: Pixel = 108;
			1829: Pixel = 112;
			1830: Pixel = 113;
			1831: Pixel = 117;
			1832: Pixel = 116;
			1833: Pixel = 112;
			1834: Pixel = 113;
			1835: Pixel = 124;
			1836: Pixel = 128;
			1837: Pixel = 131;
			1838: Pixel = 137;
			1839: Pixel = 140;
			1840: Pixel = 145;
			1841: Pixel = 142;
			1842: Pixel = 139;
			1843: Pixel = 145;
			1844: Pixel = 162;
			1845: Pixel = 169;
			1846: Pixel = 156;
			1847: Pixel = 175;
			1848: Pixel = 203;
			1849: Pixel = 205;
			1850: Pixel = 203;
			1851: Pixel = 205;
			1852: Pixel = 202;
			1853: Pixel = 199;
			1854: Pixel = 202;
			1855: Pixel = 206;
			1856: Pixel = 209;
			1857: Pixel = 210;
			1858: Pixel = 215;
			1859: Pixel = 227;
			1860: Pixel = 134;
			1861: Pixel = 69;
			1862: Pixel = 83;
			1863: Pixel = 89;
			1864: Pixel = 99;
			1865: Pixel = 129;
			1866: Pixel = 149;
			1867: Pixel = 155;
			1868: Pixel = 153;
			1869: Pixel = 153;
			1870: Pixel = 144;
			1871: Pixel = 106;
			1872: Pixel = 44;
			1873: Pixel = 59;
			1874: Pixel = 110;
			1875: Pixel = 138;
			1876: Pixel = 148;
			1877: Pixel = 144;
			1878: Pixel = 142;
			1879: Pixel = 143;
			1880: Pixel = 144;
			1881: Pixel = 144;
			1882: Pixel = 157;
			1883: Pixel = 124;
			1884: Pixel = 39;
			1885: Pixel = 45;
			1886: Pixel = 50;
			1887: Pixel = 54;
			1888: Pixel = 53;
			1889: Pixel = 44;
			1890: Pixel = 49;
			1891: Pixel = 54;
			1892: Pixel = 48;
			1893: Pixel = 53;
			1894: Pixel = 59;
			1895: Pixel = 82;
			1896: Pixel = 128;
			1897: Pixel = 150;
			1898: Pixel = 142;
			1899: Pixel = 154;
			1900: Pixel = 86;
			1901: Pixel = 88;
			1902: Pixel = 92;
			1903: Pixel = 89;
			1904: Pixel = 89;
			1905: Pixel = 121;
			1906: Pixel = 151;
			1907: Pixel = 163;
			1908: Pixel = 166;
			1909: Pixel = 165;
			1910: Pixel = 155;
			1911: Pixel = 131;
			1912: Pixel = 94;
			1913: Pixel = 75;
			1914: Pixel = 90;
			1915: Pixel = 97;
			1916: Pixel = 100;
			1917: Pixel = 99;
			1918: Pixel = 100;
			1919: Pixel = 102;
			1920: Pixel = 104;
			1921: Pixel = 109;
			1922: Pixel = 115;
			1923: Pixel = 117;
			1924: Pixel = 118;
			1925: Pixel = 120;
			1926: Pixel = 127;
			1927: Pixel = 111;
			1928: Pixel = 113;
			1929: Pixel = 112;
			1930: Pixel = 112;
			1931: Pixel = 116;
			1932: Pixel = 116;
			1933: Pixel = 118;
			1934: Pixel = 122;
			1935: Pixel = 128;
			1936: Pixel = 129;
			1937: Pixel = 137;
			1938: Pixel = 137;
			1939: Pixel = 139;
			1940: Pixel = 140;
			1941: Pixel = 135;
			1942: Pixel = 139;
			1943: Pixel = 145;
			1944: Pixel = 152;
			1945: Pixel = 153;
			1946: Pixel = 181;
			1947: Pixel = 200;
			1948: Pixel = 200;
			1949: Pixel = 202;
			1950: Pixel = 200;
			1951: Pixel = 198;
			1952: Pixel = 195;
			1953: Pixel = 201;
			1954: Pixel = 202;
			1955: Pixel = 203;
			1956: Pixel = 204;
			1957: Pixel = 208;
			1958: Pixel = 208;
			1959: Pixel = 213;
			1960: Pixel = 225;
			1961: Pixel = 168;
			1962: Pixel = 73;
			1963: Pixel = 78;
			1964: Pixel = 96;
			1965: Pixel = 128;
			1966: Pixel = 149;
			1967: Pixel = 155;
			1968: Pixel = 153;
			1969: Pixel = 154;
			1970: Pixel = 145;
			1971: Pixel = 104;
			1972: Pixel = 50;
			1973: Pixel = 43;
			1974: Pixel = 76;
			1975: Pixel = 122;
			1976: Pixel = 144;
			1977: Pixel = 148;
			1978: Pixel = 142;
			1979: Pixel = 142;
			1980: Pixel = 145;
			1981: Pixel = 151;
			1982: Pixel = 148;
			1983: Pixel = 60;
			1984: Pixel = 35;
			1985: Pixel = 45;
			1986: Pixel = 56;
			1987: Pixel = 56;
			1988: Pixel = 49;
			1989: Pixel = 45;
			1990: Pixel = 56;
			1991: Pixel = 47;
			1992: Pixel = 53;
			1993: Pixel = 55;
			1994: Pixel = 65;
			1995: Pixel = 120;
			1996: Pixel = 149;
			1997: Pixel = 144;
			1998: Pixel = 154;
			1999: Pixel = 165;
			2000: Pixel = 87;
			2001: Pixel = 92;
			2002: Pixel = 92;
			2003: Pixel = 90;
			2004: Pixel = 91;
			2005: Pixel = 123;
			2006: Pixel = 151;
			2007: Pixel = 163;
			2008: Pixel = 165;
			2009: Pixel = 164;
			2010: Pixel = 156;
			2011: Pixel = 132;
			2012: Pixel = 94;
			2013: Pixel = 75;
			2014: Pixel = 89;
			2015: Pixel = 95;
			2016: Pixel = 98;
			2017: Pixel = 101;
			2018: Pixel = 99;
			2019: Pixel = 100;
			2020: Pixel = 103;
			2021: Pixel = 109;
			2022: Pixel = 114;
			2023: Pixel = 118;
			2024: Pixel = 114;
			2025: Pixel = 131;
			2026: Pixel = 123;
			2027: Pixel = 100;
			2028: Pixel = 109;
			2029: Pixel = 115;
			2030: Pixel = 112;
			2031: Pixel = 113;
			2032: Pixel = 114;
			2033: Pixel = 119;
			2034: Pixel = 127;
			2035: Pixel = 132;
			2036: Pixel = 141;
			2037: Pixel = 139;
			2038: Pixel = 139;
			2039: Pixel = 140;
			2040: Pixel = 136;
			2041: Pixel = 133;
			2042: Pixel = 132;
			2043: Pixel = 133;
			2044: Pixel = 155;
			2045: Pixel = 188;
			2046: Pixel = 201;
			2047: Pixel = 192;
			2048: Pixel = 192;
			2049: Pixel = 191;
			2050: Pixel = 192;
			2051: Pixel = 199;
			2052: Pixel = 202;
			2053: Pixel = 203;
			2054: Pixel = 205;
			2055: Pixel = 206;
			2056: Pixel = 208;
			2057: Pixel = 207;
			2058: Pixel = 207;
			2059: Pixel = 208;
			2060: Pixel = 211;
			2061: Pixel = 233;
			2062: Pixel = 149;
			2063: Pixel = 55;
			2064: Pixel = 93;
			2065: Pixel = 125;
			2066: Pixel = 148;
			2067: Pixel = 154;
			2068: Pixel = 153;
			2069: Pixel = 153;
			2070: Pixel = 143;
			2071: Pixel = 107;
			2072: Pixel = 53;
			2073: Pixel = 39;
			2074: Pixel = 46;
			2075: Pixel = 94;
			2076: Pixel = 135;
			2077: Pixel = 143;
			2078: Pixel = 137;
			2079: Pixel = 137;
			2080: Pixel = 144;
			2081: Pixel = 158;
			2082: Pixel = 93;
			2083: Pixel = 35;
			2084: Pixel = 45;
			2085: Pixel = 51;
			2086: Pixel = 54;
			2087: Pixel = 54;
			2088: Pixel = 47;
			2089: Pixel = 53;
			2090: Pixel = 48;
			2091: Pixel = 51;
			2092: Pixel = 52;
			2093: Pixel = 51;
			2094: Pixel = 111;
			2095: Pixel = 149;
			2096: Pixel = 137;
			2097: Pixel = 150;
			2098: Pixel = 166;
			2099: Pixel = 164;
			2100: Pixel = 90;
			2101: Pixel = 92;
			2102: Pixel = 92;
			2103: Pixel = 89;
			2104: Pixel = 89;
			2105: Pixel = 123;
			2106: Pixel = 151;
			2107: Pixel = 162;
			2108: Pixel = 164;
			2109: Pixel = 163;
			2110: Pixel = 158;
			2111: Pixel = 133;
			2112: Pixel = 93;
			2113: Pixel = 77;
			2114: Pixel = 88;
			2115: Pixel = 95;
			2116: Pixel = 97;
			2117: Pixel = 101;
			2118: Pixel = 101;
			2119: Pixel = 101;
			2120: Pixel = 105;
			2121: Pixel = 110;
			2122: Pixel = 114;
			2123: Pixel = 116;
			2124: Pixel = 108;
			2125: Pixel = 160;
			2126: Pixel = 113;
			2127: Pixel = 102;
			2128: Pixel = 109;
			2129: Pixel = 111;
			2130: Pixel = 113;
			2131: Pixel = 116;
			2132: Pixel = 118;
			2133: Pixel = 124;
			2134: Pixel = 126;
			2135: Pixel = 137;
			2136: Pixel = 138;
			2137: Pixel = 131;
			2138: Pixel = 138;
			2139: Pixel = 140;
			2140: Pixel = 132;
			2141: Pixel = 116;
			2142: Pixel = 128;
			2143: Pixel = 167;
			2144: Pixel = 194;
			2145: Pixel = 187;
			2146: Pixel = 189;
			2147: Pixel = 190;
			2148: Pixel = 186;
			2149: Pixel = 191;
			2150: Pixel = 194;
			2151: Pixel = 199;
			2152: Pixel = 204;
			2153: Pixel = 204;
			2154: Pixel = 203;
			2155: Pixel = 204;
			2156: Pixel = 203;
			2157: Pixel = 203;
			2158: Pixel = 205;
			2159: Pixel = 205;
			2160: Pixel = 211;
			2161: Pixel = 217;
			2162: Pixel = 223;
			2163: Pixel = 102;
			2164: Pixel = 73;
			2165: Pixel = 124;
			2166: Pixel = 146;
			2167: Pixel = 153;
			2168: Pixel = 154;
			2169: Pixel = 154;
			2170: Pixel = 143;
			2171: Pixel = 108;
			2172: Pixel = 55;
			2173: Pixel = 44;
			2174: Pixel = 42;
			2175: Pixel = 52;
			2176: Pixel = 93;
			2177: Pixel = 148;
			2178: Pixel = 166;
			2179: Pixel = 145;
			2180: Pixel = 154;
			2181: Pixel = 122;
			2182: Pixel = 44;
			2183: Pixel = 44;
			2184: Pixel = 50;
			2185: Pixel = 53;
			2186: Pixel = 54;
			2187: Pixel = 52;
			2188: Pixel = 51;
			2189: Pixel = 51;
			2190: Pixel = 51;
			2191: Pixel = 55;
			2192: Pixel = 38;
			2193: Pixel = 91;
			2194: Pixel = 151;
			2195: Pixel = 139;
			2196: Pixel = 144;
			2197: Pixel = 162;
			2198: Pixel = 161;
			2199: Pixel = 161;
			2200: Pixel = 91;
			2201: Pixel = 90;
			2202: Pixel = 89;
			2203: Pixel = 87;
			2204: Pixel = 85;
			2205: Pixel = 120;
			2206: Pixel = 151;
			2207: Pixel = 162;
			2208: Pixel = 163;
			2209: Pixel = 163;
			2210: Pixel = 158;
			2211: Pixel = 134;
			2212: Pixel = 94;
			2213: Pixel = 74;
			2214: Pixel = 88;
			2215: Pixel = 92;
			2216: Pixel = 95;
			2217: Pixel = 98;
			2218: Pixel = 98;
			2219: Pixel = 102;
			2220: Pixel = 106;
			2221: Pixel = 107;
			2222: Pixel = 113;
			2223: Pixel = 106;
			2224: Pixel = 124;
			2225: Pixel = 173;
			2226: Pixel = 100;
			2227: Pixel = 104;
			2228: Pixel = 108;
			2229: Pixel = 113;
			2230: Pixel = 111;
			2231: Pixel = 115;
			2232: Pixel = 120;
			2233: Pixel = 127;
			2234: Pixel = 135;
			2235: Pixel = 137;
			2236: Pixel = 134;
			2237: Pixel = 133;
			2238: Pixel = 137;
			2239: Pixel = 123;
			2240: Pixel = 115;
			2241: Pixel = 134;
			2242: Pixel = 178;
			2243: Pixel = 191;
			2244: Pixel = 179;
			2245: Pixel = 187;
			2246: Pixel = 183;
			2247: Pixel = 179;
			2248: Pixel = 189;
			2249: Pixel = 198;
			2250: Pixel = 197;
			2251: Pixel = 196;
			2252: Pixel = 201;
			2253: Pixel = 202;
			2254: Pixel = 198;
			2255: Pixel = 201;
			2256: Pixel = 202;
			2257: Pixel = 201;
			2258: Pixel = 207;
			2259: Pixel = 207;
			2260: Pixel = 208;
			2261: Pixel = 210;
			2262: Pixel = 233;
			2263: Pixel = 179;
			2264: Pixel = 63;
			2265: Pixel = 122;
			2266: Pixel = 146;
			2267: Pixel = 152;
			2268: Pixel = 153;
			2269: Pixel = 154;
			2270: Pixel = 145;
			2271: Pixel = 108;
			2272: Pixel = 56;
			2273: Pixel = 46;
			2274: Pixel = 35;
			2275: Pixel = 37;
			2276: Pixel = 151;
			2277: Pixel = 209;
			2278: Pixel = 206;
			2279: Pixel = 209;
			2280: Pixel = 211;
			2281: Pixel = 77;
			2282: Pixel = 36;
			2283: Pixel = 50;
			2284: Pixel = 54;
			2285: Pixel = 55;
			2286: Pixel = 55;
			2287: Pixel = 54;
			2288: Pixel = 52;
			2289: Pixel = 49;
			2290: Pixel = 57;
			2291: Pixel = 40;
			2292: Pixel = 70;
			2293: Pixel = 144;
			2294: Pixel = 144;
			2295: Pixel = 142;
			2296: Pixel = 162;
			2297: Pixel = 161;
			2298: Pixel = 158;
			2299: Pixel = 158;
			2300: Pixel = 88;
			2301: Pixel = 89;
			2302: Pixel = 91;
			2303: Pixel = 90;
			2304: Pixel = 86;
			2305: Pixel = 118;
			2306: Pixel = 150;
			2307: Pixel = 163;
			2308: Pixel = 164;
			2309: Pixel = 163;
			2310: Pixel = 157;
			2311: Pixel = 132;
			2312: Pixel = 89;
			2313: Pixel = 70;
			2314: Pixel = 83;
			2315: Pixel = 92;
			2316: Pixel = 97;
			2317: Pixel = 97;
			2318: Pixel = 97;
			2319: Pixel = 99;
			2320: Pixel = 103;
			2321: Pixel = 105;
			2322: Pixel = 112;
			2323: Pixel = 98;
			2324: Pixel = 154;
			2325: Pixel = 170;
			2326: Pixel = 96;
			2327: Pixel = 104;
			2328: Pixel = 109;
			2329: Pixel = 114;
			2330: Pixel = 115;
			2331: Pixel = 116;
			2332: Pixel = 123;
			2333: Pixel = 130;
			2334: Pixel = 129;
			2335: Pixel = 125;
			2336: Pixel = 131;
			2337: Pixel = 135;
			2338: Pixel = 121;
			2339: Pixel = 109;
			2340: Pixel = 149;
			2341: Pixel = 182;
			2342: Pixel = 175;
			2343: Pixel = 176;
			2344: Pixel = 175;
			2345: Pixel = 174;
			2346: Pixel = 182;
			2347: Pixel = 187;
			2348: Pixel = 189;
			2349: Pixel = 193;
			2350: Pixel = 195;
			2351: Pixel = 194;
			2352: Pixel = 190;
			2353: Pixel = 194;
			2354: Pixel = 198;
			2355: Pixel = 203;
			2356: Pixel = 204;
			2357: Pixel = 202;
			2358: Pixel = 200;
			2359: Pixel = 206;
			2360: Pixel = 206;
			2361: Pixel = 205;
			2362: Pixel = 214;
			2363: Pixel = 222;
			2364: Pixel = 100;
			2365: Pixel = 105;
			2366: Pixel = 149;
			2367: Pixel = 154;
			2368: Pixel = 154;
			2369: Pixel = 154;
			2370: Pixel = 144;
			2371: Pixel = 106;
			2372: Pixel = 54;
			2373: Pixel = 27;
			2374: Pixel = 58;
			2375: Pixel = 173;
			2376: Pixel = 206;
			2377: Pixel = 201;
			2378: Pixel = 217;
			2379: Pixel = 223;
			2380: Pixel = 242;
			2381: Pixel = 132;
			2382: Pixel = 31;
			2383: Pixel = 50;
			2384: Pixel = 54;
			2385: Pixel = 54;
			2386: Pixel = 51;
			2387: Pixel = 51;
			2388: Pixel = 49;
			2389: Pixel = 54;
			2390: Pixel = 51;
			2391: Pixel = 51;
			2392: Pixel = 129;
			2393: Pixel = 151;
			2394: Pixel = 140;
			2395: Pixel = 158;
			2396: Pixel = 163;
			2397: Pixel = 159;
			2398: Pixel = 158;
			2399: Pixel = 157;
			2400: Pixel = 91;
			2401: Pixel = 92;
			2402: Pixel = 95;
			2403: Pixel = 95;
			2404: Pixel = 90;
			2405: Pixel = 118;
			2406: Pixel = 149;
			2407: Pixel = 164;
			2408: Pixel = 167;
			2409: Pixel = 165;
			2410: Pixel = 157;
			2411: Pixel = 132;
			2412: Pixel = 89;
			2413: Pixel = 72;
			2414: Pixel = 82;
			2415: Pixel = 95;
			2416: Pixel = 98;
			2417: Pixel = 100;
			2418: Pixel = 100;
			2419: Pixel = 100;
			2420: Pixel = 103;
			2421: Pixel = 107;
			2422: Pixel = 114;
			2423: Pixel = 103;
			2424: Pixel = 180;
			2425: Pixel = 157;
			2426: Pixel = 93;
			2427: Pixel = 104;
			2428: Pixel = 109;
			2429: Pixel = 109;
			2430: Pixel = 113;
			2431: Pixel = 121;
			2432: Pixel = 129;
			2433: Pixel = 122;
			2434: Pixel = 119;
			2435: Pixel = 127;
			2436: Pixel = 132;
			2437: Pixel = 118;
			2438: Pixel = 113;
			2439: Pixel = 159;
			2440: Pixel = 180;
			2441: Pixel = 169;
			2442: Pixel = 165;
			2443: Pixel = 171;
			2444: Pixel = 177;
			2445: Pixel = 180;
			2446: Pixel = 179;
			2447: Pixel = 190;
			2448: Pixel = 188;
			2449: Pixel = 188;
			2450: Pixel = 188;
			2451: Pixel = 187;
			2452: Pixel = 193;
			2453: Pixel = 197;
			2454: Pixel = 197;
			2455: Pixel = 197;
			2456: Pixel = 200;
			2457: Pixel = 199;
			2458: Pixel = 203;
			2459: Pixel = 204;
			2460: Pixel = 204;
			2461: Pixel = 205;
			2462: Pixel = 205;
			2463: Pixel = 223;
			2464: Pixel = 181;
			2465: Pixel = 98;
			2466: Pixel = 145;
			2467: Pixel = 156;
			2468: Pixel = 156;
			2469: Pixel = 155;
			2470: Pixel = 143;
			2471: Pixel = 94;
			2472: Pixel = 27;
			2473: Pixel = 87;
			2474: Pixel = 195;
			2475: Pixel = 191;
			2476: Pixel = 198;
			2477: Pixel = 218;
			2478: Pixel = 212;
			2479: Pixel = 206;
			2480: Pixel = 230;
			2481: Pixel = 176;
			2482: Pixel = 33;
			2483: Pixel = 49;
			2484: Pixel = 53;
			2485: Pixel = 50;
			2486: Pixel = 48;
			2487: Pixel = 45;
			2488: Pixel = 48;
			2489: Pixel = 56;
			2490: Pixel = 45;
			2491: Pixel = 102;
			2492: Pixel = 156;
			2493: Pixel = 141;
			2494: Pixel = 154;
			2495: Pixel = 160;
			2496: Pixel = 158;
			2497: Pixel = 159;
			2498: Pixel = 157;
			2499: Pixel = 158;
			2500: Pixel = 95;
			2501: Pixel = 96;
			2502: Pixel = 98;
			2503: Pixel = 97;
			2504: Pixel = 94;
			2505: Pixel = 118;
			2506: Pixel = 149;
			2507: Pixel = 165;
			2508: Pixel = 167;
			2509: Pixel = 167;
			2510: Pixel = 160;
			2511: Pixel = 135;
			2512: Pixel = 92;
			2513: Pixel = 76;
			2514: Pixel = 88;
			2515: Pixel = 96;
			2516: Pixel = 99;
			2517: Pixel = 101;
			2518: Pixel = 101;
			2519: Pixel = 102;
			2520: Pixel = 106;
			2521: Pixel = 110;
			2522: Pixel = 112;
			2523: Pixel = 108;
			2524: Pixel = 194;
			2525: Pixel = 145;
			2526: Pixel = 94;
			2527: Pixel = 104;
			2528: Pixel = 102;
			2529: Pixel = 110;
			2530: Pixel = 119;
			2531: Pixel = 123;
			2532: Pixel = 120;
			2533: Pixel = 119;
			2534: Pixel = 130;
			2535: Pixel = 135;
			2536: Pixel = 119;
			2537: Pixel = 115;
			2538: Pixel = 157;
			2539: Pixel = 168;
			2540: Pixel = 163;
			2541: Pixel = 163;
			2542: Pixel = 167;
			2543: Pixel = 179;
			2544: Pixel = 180;
			2545: Pixel = 178;
			2546: Pixel = 186;
			2547: Pixel = 183;
			2548: Pixel = 185;
			2549: Pixel = 176;
			2550: Pixel = 179;
			2551: Pixel = 188;
			2552: Pixel = 196;
			2553: Pixel = 197;
			2554: Pixel = 194;
			2555: Pixel = 194;
			2556: Pixel = 200;
			2557: Pixel = 198;
			2558: Pixel = 190;
			2559: Pixel = 197;
			2560: Pixel = 200;
			2561: Pixel = 202;
			2562: Pixel = 203;
			2563: Pixel = 204;
			2564: Pixel = 216;
			2565: Pixel = 172;
			2566: Pixel = 138;
			2567: Pixel = 153;
			2568: Pixel = 155;
			2569: Pixel = 153;
			2570: Pixel = 124;
			2571: Pixel = 83;
			2572: Pixel = 136;
			2573: Pixel = 204;
			2574: Pixel = 191;
			2575: Pixel = 202;
			2576: Pixel = 215;
			2577: Pixel = 205;
			2578: Pixel = 200;
			2579: Pixel = 205;
			2580: Pixel = 230;
			2581: Pixel = 175;
			2582: Pixel = 34;
			2583: Pixel = 53;
			2584: Pixel = 54;
			2585: Pixel = 46;
			2586: Pixel = 45;
			2587: Pixel = 48;
			2588: Pixel = 54;
			2589: Pixel = 38;
			2590: Pixel = 63;
			2591: Pixel = 148;
			2592: Pixel = 148;
			2593: Pixel = 150;
			2594: Pixel = 161;
			2595: Pixel = 157;
			2596: Pixel = 157;
			2597: Pixel = 157;
			2598: Pixel = 155;
			2599: Pixel = 156;
			2600: Pixel = 98;
			2601: Pixel = 100;
			2602: Pixel = 100;
			2603: Pixel = 98;
			2604: Pixel = 95;
			2605: Pixel = 119;
			2606: Pixel = 149;
			2607: Pixel = 163;
			2608: Pixel = 167;
			2609: Pixel = 168;
			2610: Pixel = 163;
			2611: Pixel = 136;
			2612: Pixel = 93;
			2613: Pixel = 77;
			2614: Pixel = 88;
			2615: Pixel = 97;
			2616: Pixel = 101;
			2617: Pixel = 102;
			2618: Pixel = 103;
			2619: Pixel = 99;
			2620: Pixel = 106;
			2621: Pixel = 111;
			2622: Pixel = 108;
			2623: Pixel = 119;
			2624: Pixel = 197;
			2625: Pixel = 128;
			2626: Pixel = 97;
			2627: Pixel = 100;
			2628: Pixel = 107;
			2629: Pixel = 109;
			2630: Pixel = 113;
			2631: Pixel = 116;
			2632: Pixel = 122;
			2633: Pixel = 127;
			2634: Pixel = 124;
			2635: Pixel = 115;
			2636: Pixel = 117;
			2637: Pixel = 156;
			2638: Pixel = 157;
			2639: Pixel = 148;
			2640: Pixel = 151;
			2641: Pixel = 164;
			2642: Pixel = 173;
			2643: Pixel = 177;
			2644: Pixel = 179;
			2645: Pixel = 177;
			2646: Pixel = 179;
			2647: Pixel = 181;
			2648: Pixel = 169;
			2649: Pixel = 177;
			2650: Pixel = 185;
			2651: Pixel = 186;
			2652: Pixel = 186;
			2653: Pixel = 192;
			2654: Pixel = 194;
			2655: Pixel = 201;
			2656: Pixel = 197;
			2657: Pixel = 176;
			2658: Pixel = 182;
			2659: Pixel = 199;
			2660: Pixel = 200;
			2661: Pixel = 201;
			2662: Pixel = 200;
			2663: Pixel = 197;
			2664: Pixel = 200;
			2665: Pixel = 218;
			2666: Pixel = 175;
			2667: Pixel = 148;
			2668: Pixel = 149;
			2669: Pixel = 142;
			2670: Pixel = 152;
			2671: Pixel = 189;
			2672: Pixel = 204;
			2673: Pixel = 192;
			2674: Pixel = 209;
			2675: Pixel = 209;
			2676: Pixel = 201;
			2677: Pixel = 201;
			2678: Pixel = 205;
			2679: Pixel = 211;
			2680: Pixel = 233;
			2681: Pixel = 153;
			2682: Pixel = 33;
			2683: Pixel = 51;
			2684: Pixel = 52;
			2685: Pixel = 51;
			2686: Pixel = 44;
			2687: Pixel = 52;
			2688: Pixel = 50;
			2689: Pixel = 36;
			2690: Pixel = 118;
			2691: Pixel = 156;
			2692: Pixel = 146;
			2693: Pixel = 160;
			2694: Pixel = 159;
			2695: Pixel = 157;
			2696: Pixel = 156;
			2697: Pixel = 156;
			2698: Pixel = 155;
			2699: Pixel = 154;
			2700: Pixel = 99;
			2701: Pixel = 99;
			2702: Pixel = 99;
			2703: Pixel = 98;
			2704: Pixel = 98;
			2705: Pixel = 123;
			2706: Pixel = 150;
			2707: Pixel = 163;
			2708: Pixel = 169;
			2709: Pixel = 171;
			2710: Pixel = 165;
			2711: Pixel = 138;
			2712: Pixel = 93;
			2713: Pixel = 77;
			2714: Pixel = 90;
			2715: Pixel = 97;
			2716: Pixel = 100;
			2717: Pixel = 101;
			2718: Pixel = 100;
			2719: Pixel = 99;
			2720: Pixel = 103;
			2721: Pixel = 109;
			2722: Pixel = 97;
			2723: Pixel = 132;
			2724: Pixel = 192;
			2725: Pixel = 127;
			2726: Pixel = 106;
			2727: Pixel = 104;
			2728: Pixel = 103;
			2729: Pixel = 102;
			2730: Pixel = 109;
			2731: Pixel = 115;
			2732: Pixel = 121;
			2733: Pixel = 120;
			2734: Pixel = 115;
			2735: Pixel = 125;
			2736: Pixel = 149;
			2737: Pixel = 152;
			2738: Pixel = 147;
			2739: Pixel = 143;
			2740: Pixel = 153;
			2741: Pixel = 165;
			2742: Pixel = 175;
			2743: Pixel = 171;
			2744: Pixel = 165;
			2745: Pixel = 178;
			2746: Pixel = 176;
			2747: Pixel = 165;
			2748: Pixel = 176;
			2749: Pixel = 178;
			2750: Pixel = 181;
			2751: Pixel = 178;
			2752: Pixel = 178;
			2753: Pixel = 184;
			2754: Pixel = 188;
			2755: Pixel = 186;
			2756: Pixel = 181;
			2757: Pixel = 182;
			2758: Pixel = 188;
			2759: Pixel = 192;
			2760: Pixel = 196;
			2761: Pixel = 195;
			2762: Pixel = 193;
			2763: Pixel = 195;
			2764: Pixel = 189;
			2765: Pixel = 195;
			2766: Pixel = 194;
			2767: Pixel = 148;
			2768: Pixel = 156;
			2769: Pixel = 185;
			2770: Pixel = 203;
			2771: Pixel = 193;
			2772: Pixel = 197;
			2773: Pixel = 208;
			2774: Pixel = 203;
			2775: Pixel = 200;
			2776: Pixel = 202;
			2777: Pixel = 203;
			2778: Pixel = 207;
			2779: Pixel = 213;
			2780: Pixel = 233;
			2781: Pixel = 123;
			2782: Pixel = 36;
			2783: Pixel = 55;
			2784: Pixel = 50;
			2785: Pixel = 46;
			2786: Pixel = 44;
			2787: Pixel = 51;
			2788: Pixel = 49;
			2789: Pixel = 86;
			2790: Pixel = 151;
			2791: Pixel = 146;
			2792: Pixel = 154;
			2793: Pixel = 161;
			2794: Pixel = 158;
			2795: Pixel = 157;
			2796: Pixel = 157;
			2797: Pixel = 155;
			2798: Pixel = 154;
			2799: Pixel = 153;
			2800: Pixel = 100;
			2801: Pixel = 100;
			2802: Pixel = 98;
			2803: Pixel = 99;
			2804: Pixel = 100;
			2805: Pixel = 123;
			2806: Pixel = 152;
			2807: Pixel = 167;
			2808: Pixel = 172;
			2809: Pixel = 173;
			2810: Pixel = 168;
			2811: Pixel = 140;
			2812: Pixel = 93;
			2813: Pixel = 76;
			2814: Pixel = 90;
			2815: Pixel = 95;
			2816: Pixel = 99;
			2817: Pixel = 100;
			2818: Pixel = 98;
			2819: Pixel = 99;
			2820: Pixel = 101;
			2821: Pixel = 107;
			2822: Pixel = 90;
			2823: Pixel = 153;
			2824: Pixel = 197;
			2825: Pixel = 136;
			2826: Pixel = 109;
			2827: Pixel = 105;
			2828: Pixel = 105;
			2829: Pixel = 108;
			2830: Pixel = 113;
			2831: Pixel = 117;
			2832: Pixel = 121;
			2833: Pixel = 119;
			2834: Pixel = 123;
			2835: Pixel = 150;
			2836: Pixel = 148;
			2837: Pixel = 140;
			2838: Pixel = 137;
			2839: Pixel = 145;
			2840: Pixel = 162;
			2841: Pixel = 161;
			2842: Pixel = 159;
			2843: Pixel = 171;
			2844: Pixel = 176;
			2845: Pixel = 162;
			2846: Pixel = 165;
			2847: Pixel = 174;
			2848: Pixel = 175;
			2849: Pixel = 175;
			2850: Pixel = 173;
			2851: Pixel = 175;
			2852: Pixel = 183;
			2853: Pixel = 187;
			2854: Pixel = 177;
			2855: Pixel = 177;
			2856: Pixel = 187;
			2857: Pixel = 184;
			2858: Pixel = 189;
			2859: Pixel = 192;
			2860: Pixel = 189;
			2861: Pixel = 184;
			2862: Pixel = 186;
			2863: Pixel = 188;
			2864: Pixel = 184;
			2865: Pixel = 180;
			2866: Pixel = 190;
			2867: Pixel = 184;
			2868: Pixel = 197;
			2869: Pixel = 195;
			2870: Pixel = 196;
			2871: Pixel = 204;
			2872: Pixel = 206;
			2873: Pixel = 200;
			2874: Pixel = 199;
			2875: Pixel = 202;
			2876: Pixel = 205;
			2877: Pixel = 201;
			2878: Pixel = 203;
			2879: Pixel = 213;
			2880: Pixel = 230;
			2881: Pixel = 91;
			2882: Pixel = 37;
			2883: Pixel = 53;
			2884: Pixel = 52;
			2885: Pixel = 44;
			2886: Pixel = 49;
			2887: Pixel = 54;
			2888: Pixel = 72;
			2889: Pixel = 134;
			2890: Pixel = 149;
			2891: Pixel = 148;
			2892: Pixel = 160;
			2893: Pixel = 159;
			2894: Pixel = 158;
			2895: Pixel = 156;
			2896: Pixel = 156;
			2897: Pixel = 154;
			2898: Pixel = 154;
			2899: Pixel = 154;
			2900: Pixel = 98;
			2901: Pixel = 99;
			2902: Pixel = 97;
			2903: Pixel = 97;
			2904: Pixel = 99;
			2905: Pixel = 120;
			2906: Pixel = 150;
			2907: Pixel = 168;
			2908: Pixel = 173;
			2909: Pixel = 174;
			2910: Pixel = 167;
			2911: Pixel = 138;
			2912: Pixel = 94;
			2913: Pixel = 75;
			2914: Pixel = 88;
			2915: Pixel = 95;
			2916: Pixel = 98;
			2917: Pixel = 98;
			2918: Pixel = 98;
			2919: Pixel = 98;
			2920: Pixel = 101;
			2921: Pixel = 107;
			2922: Pixel = 89;
			2923: Pixel = 169;
			2924: Pixel = 194;
			2925: Pixel = 143;
			2926: Pixel = 126;
			2927: Pixel = 114;
			2928: Pixel = 104;
			2929: Pixel = 109;
			2930: Pixel = 109;
			2931: Pixel = 119;
			2932: Pixel = 118;
			2933: Pixel = 120;
			2934: Pixel = 145;
			2935: Pixel = 144;
			2936: Pixel = 141;
			2937: Pixel = 133;
			2938: Pixel = 145;
			2939: Pixel = 152;
			2940: Pixel = 145;
			2941: Pixel = 151;
			2942: Pixel = 171;
			2943: Pixel = 170;
			2944: Pixel = 159;
			2945: Pixel = 168;
			2946: Pixel = 171;
			2947: Pixel = 171;
			2948: Pixel = 175;
			2949: Pixel = 174;
			2950: Pixel = 173;
			2951: Pixel = 169;
			2952: Pixel = 176;
			2953: Pixel = 181;
			2954: Pixel = 181;
			2955: Pixel = 182;
			2956: Pixel = 180;
			2957: Pixel = 190;
			2958: Pixel = 187;
			2959: Pixel = 184;
			2960: Pixel = 177;
			2961: Pixel = 175;
			2962: Pixel = 185;
			2963: Pixel = 175;
			2964: Pixel = 167;
			2965: Pixel = 179;
			2966: Pixel = 189;
			2967: Pixel = 189;
			2968: Pixel = 196;
			2969: Pixel = 204;
			2970: Pixel = 207;
			2971: Pixel = 197;
			2972: Pixel = 199;
			2973: Pixel = 198;
			2974: Pixel = 200;
			2975: Pixel = 205;
			2976: Pixel = 200;
			2977: Pixel = 178;
			2978: Pixel = 202;
			2979: Pixel = 215;
			2980: Pixel = 206;
			2981: Pixel = 54;
			2982: Pixel = 39;
			2983: Pixel = 50;
			2984: Pixel = 51;
			2985: Pixel = 45;
			2986: Pixel = 54;
			2987: Pixel = 45;
			2988: Pixel = 105;
			2989: Pixel = 154;
			2990: Pixel = 145;
			2991: Pixel = 157;
			2992: Pixel = 161;
			2993: Pixel = 159;
			2994: Pixel = 159;
			2995: Pixel = 157;
			2996: Pixel = 158;
			2997: Pixel = 157;
			2998: Pixel = 156;
			2999: Pixel = 157;
			3000: Pixel = 97;
			3001: Pixel = 97;
			3002: Pixel = 97;
			3003: Pixel = 97;
			3004: Pixel = 97;
			3005: Pixel = 121;
			3006: Pixel = 152;
			3007: Pixel = 169;
			3008: Pixel = 172;
			3009: Pixel = 172;
			3010: Pixel = 166;
			3011: Pixel = 140;
			3012: Pixel = 95;
			3013: Pixel = 78;
			3014: Pixel = 92;
			3015: Pixel = 96;
			3016: Pixel = 100;
			3017: Pixel = 99;
			3018: Pixel = 98;
			3019: Pixel = 98;
			3020: Pixel = 101;
			3021: Pixel = 105;
			3022: Pixel = 90;
			3023: Pixel = 170;
			3024: Pixel = 190;
			3025: Pixel = 153;
			3026: Pixel = 140;
			3027: Pixel = 125;
			3028: Pixel = 106;
			3029: Pixel = 99;
			3030: Pixel = 114;
			3031: Pixel = 112;
			3032: Pixel = 116;
			3033: Pixel = 142;
			3034: Pixel = 141;
			3035: Pixel = 140;
			3036: Pixel = 125;
			3037: Pixel = 144;
			3038: Pixel = 151;
			3039: Pixel = 149;
			3040: Pixel = 145;
			3041: Pixel = 149;
			3042: Pixel = 157;
			3043: Pixel = 156;
			3044: Pixel = 168;
			3045: Pixel = 172;
			3046: Pixel = 166;
			3047: Pixel = 167;
			3048: Pixel = 172;
			3049: Pixel = 169;
			3050: Pixel = 165;
			3051: Pixel = 168;
			3052: Pixel = 165;
			3053: Pixel = 169;
			3054: Pixel = 172;
			3055: Pixel = 179;
			3056: Pixel = 183;
			3057: Pixel = 182;
			3058: Pixel = 179;
			3059: Pixel = 173;
			3060: Pixel = 184;
			3061: Pixel = 171;
			3062: Pixel = 166;
			3063: Pixel = 171;
			3064: Pixel = 183;
			3065: Pixel = 190;
			3066: Pixel = 191;
			3067: Pixel = 199;
			3068: Pixel = 202;
			3069: Pixel = 198;
			3070: Pixel = 195;
			3071: Pixel = 198;
			3072: Pixel = 199;
			3073: Pixel = 200;
			3074: Pixel = 203;
			3075: Pixel = 207;
			3076: Pixel = 172;
			3077: Pixel = 163;
			3078: Pixel = 171;
			3079: Pixel = 204;
			3080: Pixel = 152;
			3081: Pixel = 35;
			3082: Pixel = 51;
			3083: Pixel = 51;
			3084: Pixel = 47;
			3085: Pixel = 46;
			3086: Pixel = 50;
			3087: Pixel = 71;
			3088: Pixel = 140;
			3089: Pixel = 149;
			3090: Pixel = 151;
			3091: Pixel = 161;
			3092: Pixel = 160;
			3093: Pixel = 160;
			3094: Pixel = 159;
			3095: Pixel = 157;
			3096: Pixel = 157;
			3097: Pixel = 158;
			3098: Pixel = 157;
			3099: Pixel = 156;
			3100: Pixel = 97;
			3101: Pixel = 94;
			3102: Pixel = 94;
			3103: Pixel = 95;
			3104: Pixel = 97;
			3105: Pixel = 123;
			3106: Pixel = 154;
			3107: Pixel = 168;
			3108: Pixel = 170;
			3109: Pixel = 171;
			3110: Pixel = 166;
			3111: Pixel = 140;
			3112: Pixel = 94;
			3113: Pixel = 77;
			3114: Pixel = 91;
			3115: Pixel = 98;
			3116: Pixel = 99;
			3117: Pixel = 98;
			3118: Pixel = 98;
			3119: Pixel = 98;
			3120: Pixel = 101;
			3121: Pixel = 101;
			3122: Pixel = 87;
			3123: Pixel = 171;
			3124: Pixel = 185;
			3125: Pixel = 157;
			3126: Pixel = 144;
			3127: Pixel = 134;
			3128: Pixel = 107;
			3129: Pixel = 100;
			3130: Pixel = 106;
			3131: Pixel = 119;
			3132: Pixel = 141;
			3133: Pixel = 135;
			3134: Pixel = 135;
			3135: Pixel = 123;
			3136: Pixel = 137;
			3137: Pixel = 148;
			3138: Pixel = 143;
			3139: Pixel = 141;
			3140: Pixel = 151;
			3141: Pixel = 149;
			3142: Pixel = 145;
			3143: Pixel = 160;
			3144: Pixel = 162;
			3145: Pixel = 164;
			3146: Pixel = 167;
			3147: Pixel = 166;
			3148: Pixel = 163;
			3149: Pixel = 165;
			3150: Pixel = 160;
			3151: Pixel = 161;
			3152: Pixel = 161;
			3153: Pixel = 165;
			3154: Pixel = 173;
			3155: Pixel = 168;
			3156: Pixel = 175;
			3157: Pixel = 173;
			3158: Pixel = 171;
			3159: Pixel = 168;
			3160: Pixel = 167;
			3161: Pixel = 165;
			3162: Pixel = 173;
			3163: Pixel = 184;
			3164: Pixel = 189;
			3165: Pixel = 199;
			3166: Pixel = 204;
			3167: Pixel = 196;
			3168: Pixel = 192;
			3169: Pixel = 191;
			3170: Pixel = 196;
			3171: Pixel = 200;
			3172: Pixel = 200;
			3173: Pixel = 201;
			3174: Pixel = 210;
			3175: Pixel = 188;
			3176: Pixel = 160;
			3177: Pixel = 162;
			3178: Pixel = 147;
			3179: Pixel = 201;
			3180: Pixel = 91;
			3181: Pixel = 31;
			3182: Pixel = 56;
			3183: Pixel = 47;
			3184: Pixel = 45;
			3185: Pixel = 47;
			3186: Pixel = 59;
			3187: Pixel = 123;
			3188: Pixel = 153;
			3189: Pixel = 145;
			3190: Pixel = 158;
			3191: Pixel = 161;
			3192: Pixel = 158;
			3193: Pixel = 158;
			3194: Pixel = 158;
			3195: Pixel = 158;
			3196: Pixel = 156;
			3197: Pixel = 157;
			3198: Pixel = 157;
			3199: Pixel = 156;
			3200: Pixel = 97;
			3201: Pixel = 95;
			3202: Pixel = 95;
			3203: Pixel = 94;
			3204: Pixel = 99;
			3205: Pixel = 125;
			3206: Pixel = 153;
			3207: Pixel = 168;
			3208: Pixel = 171;
			3209: Pixel = 172;
			3210: Pixel = 166;
			3211: Pixel = 143;
			3212: Pixel = 96;
			3213: Pixel = 77;
			3214: Pixel = 91;
			3215: Pixel = 97;
			3216: Pixel = 97;
			3217: Pixel = 97;
			3218: Pixel = 97;
			3219: Pixel = 99;
			3220: Pixel = 99;
			3221: Pixel = 98;
			3222: Pixel = 87;
			3223: Pixel = 181;
			3224: Pixel = 189;
			3225: Pixel = 162;
			3226: Pixel = 147;
			3227: Pixel = 137;
			3228: Pixel = 120;
			3229: Pixel = 102;
			3230: Pixel = 115;
			3231: Pixel = 138;
			3232: Pixel = 137;
			3233: Pixel = 130;
			3234: Pixel = 119;
			3235: Pixel = 137;
			3236: Pixel = 147;
			3237: Pixel = 139;
			3238: Pixel = 132;
			3239: Pixel = 142;
			3240: Pixel = 145;
			3241: Pixel = 145;
			3242: Pixel = 162;
			3243: Pixel = 156;
			3244: Pixel = 157;
			3245: Pixel = 162;
			3246: Pixel = 151;
			3247: Pixel = 149;
			3248: Pixel = 157;
			3249: Pixel = 159;
			3250: Pixel = 156;
			3251: Pixel = 163;
			3252: Pixel = 165;
			3253: Pixel = 165;
			3254: Pixel = 164;
			3255: Pixel = 168;
			3256: Pixel = 164;
			3257: Pixel = 164;
			3258: Pixel = 162;
			3259: Pixel = 157;
			3260: Pixel = 166;
			3261: Pixel = 181;
			3262: Pixel = 184;
			3263: Pixel = 192;
			3264: Pixel = 196;
			3265: Pixel = 192;
			3266: Pixel = 189;
			3267: Pixel = 192;
			3268: Pixel = 195;
			3269: Pixel = 198;
			3270: Pixel = 202;
			3271: Pixel = 202;
			3272: Pixel = 201;
			3273: Pixel = 206;
			3274: Pixel = 206;
			3275: Pixel = 165;
			3276: Pixel = 166;
			3277: Pixel = 149;
			3278: Pixel = 159;
			3279: Pixel = 189;
			3280: Pixel = 49;
			3281: Pixel = 45;
			3282: Pixel = 50;
			3283: Pixel = 50;
			3284: Pixel = 53;
			3285: Pixel = 48;
			3286: Pixel = 84;
			3287: Pixel = 150;
			3288: Pixel = 146;
			3289: Pixel = 152;
			3290: Pixel = 160;
			3291: Pixel = 158;
			3292: Pixel = 156;
			3293: Pixel = 156;
			3294: Pixel = 158;
			3295: Pixel = 157;
			3296: Pixel = 156;
			3297: Pixel = 156;
			3298: Pixel = 156;
			3299: Pixel = 156;
			3300: Pixel = 97;
			3301: Pixel = 98;
			3302: Pixel = 96;
			3303: Pixel = 99;
			3304: Pixel = 105;
			3305: Pixel = 125;
			3306: Pixel = 153;
			3307: Pixel = 168;
			3308: Pixel = 172;
			3309: Pixel = 172;
			3310: Pixel = 167;
			3311: Pixel = 144;
			3312: Pixel = 95;
			3313: Pixel = 73;
			3314: Pixel = 89;
			3315: Pixel = 97;
			3316: Pixel = 97;
			3317: Pixel = 95;
			3318: Pixel = 97;
			3319: Pixel = 97;
			3320: Pixel = 98;
			3321: Pixel = 96;
			3322: Pixel = 85;
			3323: Pixel = 189;
			3324: Pixel = 198;
			3325: Pixel = 171;
			3326: Pixel = 157;
			3327: Pixel = 151;
			3328: Pixel = 131;
			3329: Pixel = 104;
			3330: Pixel = 132;
			3331: Pixel = 131;
			3332: Pixel = 130;
			3333: Pixel = 119;
			3334: Pixel = 137;
			3335: Pixel = 142;
			3336: Pixel = 138;
			3337: Pixel = 128;
			3338: Pixel = 135;
			3339: Pixel = 144;
			3340: Pixel = 139;
			3341: Pixel = 154;
			3342: Pixel = 139;
			3343: Pixel = 130;
			3344: Pixel = 126;
			3345: Pixel = 134;
			3346: Pixel = 134;
			3347: Pixel = 139;
			3348: Pixel = 115;
			3349: Pixel = 146;
			3350: Pixel = 163;
			3351: Pixel = 160;
			3352: Pixel = 158;
			3353: Pixel = 162;
			3354: Pixel = 165;
			3355: Pixel = 146;
			3356: Pixel = 152;
			3357: Pixel = 154;
			3358: Pixel = 153;
			3359: Pixel = 175;
			3360: Pixel = 181;
			3361: Pixel = 187;
			3362: Pixel = 197;
			3363: Pixel = 196;
			3364: Pixel = 188;
			3365: Pixel = 188;
			3366: Pixel = 193;
			3367: Pixel = 197;
			3368: Pixel = 199;
			3369: Pixel = 201;
			3370: Pixel = 203;
			3371: Pixel = 201;
			3372: Pixel = 203;
			3373: Pixel = 216;
			3374: Pixel = 190;
			3375: Pixel = 150;
			3376: Pixel = 118;
			3377: Pixel = 100;
			3378: Pixel = 188;
			3379: Pixel = 146;
			3380: Pixel = 24;
			3381: Pixel = 52;
			3382: Pixel = 49;
			3383: Pixel = 52;
			3384: Pixel = 56;
			3385: Pixel = 53;
			3386: Pixel = 121;
			3387: Pixel = 154;
			3388: Pixel = 146;
			3389: Pixel = 158;
			3390: Pixel = 159;
			3391: Pixel = 157;
			3392: Pixel = 156;
			3393: Pixel = 155;
			3394: Pixel = 156;
			3395: Pixel = 155;
			3396: Pixel = 155;
			3397: Pixel = 156;
			3398: Pixel = 155;
			3399: Pixel = 154;
			3400: Pixel = 99;
			3401: Pixel = 97;
			3402: Pixel = 98;
			3403: Pixel = 100;
			3404: Pixel = 105;
			3405: Pixel = 128;
			3406: Pixel = 154;
			3407: Pixel = 169;
			3408: Pixel = 173;
			3409: Pixel = 173;
			3410: Pixel = 169;
			3411: Pixel = 144;
			3412: Pixel = 94;
			3413: Pixel = 73;
			3414: Pixel = 87;
			3415: Pixel = 96;
			3416: Pixel = 97;
			3417: Pixel = 99;
			3418: Pixel = 99;
			3419: Pixel = 98;
			3420: Pixel = 99;
			3421: Pixel = 95;
			3422: Pixel = 83;
			3423: Pixel = 187;
			3424: Pixel = 202;
			3425: Pixel = 178;
			3426: Pixel = 155;
			3427: Pixel = 151;
			3428: Pixel = 141;
			3429: Pixel = 116;
			3430: Pixel = 122;
			3431: Pixel = 125;
			3432: Pixel = 115;
			3433: Pixel = 133;
			3434: Pixel = 141;
			3435: Pixel = 133;
			3436: Pixel = 123;
			3437: Pixel = 131;
			3438: Pixel = 137;
			3439: Pixel = 134;
			3440: Pixel = 150;
			3441: Pixel = 135;
			3442: Pixel = 124;
			3443: Pixel = 124;
			3444: Pixel = 104;
			3445: Pixel = 81;
			3446: Pixel = 96;
			3447: Pixel = 171;
			3448: Pixel = 147;
			3449: Pixel = 119;
			3450: Pixel = 111;
			3451: Pixel = 116;
			3452: Pixel = 124;
			3453: Pixel = 107;
			3454: Pixel = 98;
			3455: Pixel = 80;
			3456: Pixel = 64;
			3457: Pixel = 157;
			3458: Pixel = 170;
			3459: Pixel = 173;
			3460: Pixel = 190;
			3461: Pixel = 200;
			3462: Pixel = 194;
			3463: Pixel = 193;
			3464: Pixel = 192;
			3465: Pixel = 194;
			3466: Pixel = 198;
			3467: Pixel = 200;
			3468: Pixel = 200;
			3469: Pixel = 202;
			3470: Pixel = 204;
			3471: Pixel = 210;
			3472: Pixel = 213;
			3473: Pixel = 189;
			3474: Pixel = 131;
			3475: Pixel = 90;
			3476: Pixel = 81;
			3477: Pixel = 151;
			3478: Pixel = 213;
			3479: Pixel = 61;
			3480: Pixel = 38;
			3481: Pixel = 49;
			3482: Pixel = 44;
			3483: Pixel = 52;
			3484: Pixel = 47;
			3485: Pixel = 78;
			3486: Pixel = 148;
			3487: Pixel = 146;
			3488: Pixel = 154;
			3489: Pixel = 161;
			3490: Pixel = 158;
			3491: Pixel = 158;
			3492: Pixel = 156;
			3493: Pixel = 156;
			3494: Pixel = 155;
			3495: Pixel = 154;
			3496: Pixel = 154;
			3497: Pixel = 154;
			3498: Pixel = 153;
			3499: Pixel = 153;
			3500: Pixel = 99;
			3501: Pixel = 101;
			3502: Pixel = 98;
			3503: Pixel = 101;
			3504: Pixel = 108;
			3505: Pixel = 129;
			3506: Pixel = 156;
			3507: Pixel = 170;
			3508: Pixel = 172;
			3509: Pixel = 173;
			3510: Pixel = 169;
			3511: Pixel = 145;
			3512: Pixel = 95;
			3513: Pixel = 73;
			3514: Pixel = 87;
			3515: Pixel = 96;
			3516: Pixel = 98;
			3517: Pixel = 99;
			3518: Pixel = 99;
			3519: Pixel = 98;
			3520: Pixel = 99;
			3521: Pixel = 99;
			3522: Pixel = 81;
			3523: Pixel = 173;
			3524: Pixel = 207;
			3525: Pixel = 193;
			3526: Pixel = 149;
			3527: Pixel = 127;
			3528: Pixel = 129;
			3529: Pixel = 110;
			3530: Pixel = 121;
			3531: Pixel = 108;
			3532: Pixel = 128;
			3533: Pixel = 139;
			3534: Pixel = 131;
			3535: Pixel = 124;
			3536: Pixel = 132;
			3537: Pixel = 132;
			3538: Pixel = 129;
			3539: Pixel = 145;
			3540: Pixel = 127;
			3541: Pixel = 126;
			3542: Pixel = 133;
			3543: Pixel = 112;
			3544: Pixel = 110;
			3545: Pixel = 98;
			3546: Pixel = 87;
			3547: Pixel = 121;
			3548: Pixel = 119;
			3549: Pixel = 80;
			3550: Pixel = 78;
			3551: Pixel = 82;
			3552: Pixel = 67;
			3553: Pixel = 53;
			3554: Pixel = 32;
			3555: Pixel = 40;
			3556: Pixel = 109;
			3557: Pixel = 161;
			3558: Pixel = 179;
			3559: Pixel = 198;
			3560: Pixel = 197;
			3561: Pixel = 192;
			3562: Pixel = 194;
			3563: Pixel = 195;
			3564: Pixel = 191;
			3565: Pixel = 194;
			3566: Pixel = 198;
			3567: Pixel = 198;
			3568: Pixel = 198;
			3569: Pixel = 209;
			3570: Pixel = 206;
			3571: Pixel = 171;
			3572: Pixel = 126;
			3573: Pixel = 94;
			3574: Pixel = 81;
			3575: Pixel = 93;
			3576: Pixel = 145;
			3577: Pixel = 208;
			3578: Pixel = 113;
			3579: Pixel = 32;
			3580: Pixel = 52;
			3581: Pixel = 49;
			3582: Pixel = 48;
			3583: Pixel = 51;
			3584: Pixel = 41;
			3585: Pixel = 116;
			3586: Pixel = 151;
			3587: Pixel = 146;
			3588: Pixel = 162;
			3589: Pixel = 160;
			3590: Pixel = 159;
			3591: Pixel = 159;
			3592: Pixel = 157;
			3593: Pixel = 156;
			3594: Pixel = 154;
			3595: Pixel = 154;
			3596: Pixel = 154;
			3597: Pixel = 154;
			3598: Pixel = 153;
			3599: Pixel = 153;
			3600: Pixel = 102;
			3601: Pixel = 103;
			3602: Pixel = 97;
			3603: Pixel = 100;
			3604: Pixel = 109;
			3605: Pixel = 129;
			3606: Pixel = 154;
			3607: Pixel = 170;
			3608: Pixel = 171;
			3609: Pixel = 172;
			3610: Pixel = 169;
			3611: Pixel = 145;
			3612: Pixel = 94;
			3613: Pixel = 74;
			3614: Pixel = 89;
			3615: Pixel = 96;
			3616: Pixel = 98;
			3617: Pixel = 98;
			3618: Pixel = 100;
			3619: Pixel = 99;
			3620: Pixel = 99;
			3621: Pixel = 98;
			3622: Pixel = 79;
			3623: Pixel = 147;
			3624: Pixel = 214;
			3625: Pixel = 197;
			3626: Pixel = 147;
			3627: Pixel = 126;
			3628: Pixel = 140;
			3629: Pixel = 122;
			3630: Pixel = 106;
			3631: Pixel = 122;
			3632: Pixel = 140;
			3633: Pixel = 131;
			3634: Pixel = 121;
			3635: Pixel = 130;
			3636: Pixel = 133;
			3637: Pixel = 128;
			3638: Pixel = 138;
			3639: Pixel = 126;
			3640: Pixel = 122;
			3641: Pixel = 134;
			3642: Pixel = 108;
			3643: Pixel = 108;
			3644: Pixel = 87;
			3645: Pixel = 66;
			3646: Pixel = 61;
			3647: Pixel = 100;
			3648: Pixel = 99;
			3649: Pixel = 87;
			3650: Pixel = 102;
			3651: Pixel = 71;
			3652: Pixel = 75;
			3653: Pixel = 42;
			3654: Pixel = 42;
			3655: Pixel = 126;
			3656: Pixel = 155;
			3657: Pixel = 176;
			3658: Pixel = 192;
			3659: Pixel = 194;
			3660: Pixel = 193;
			3661: Pixel = 191;
			3662: Pixel = 191;
			3663: Pixel = 192;
			3664: Pixel = 192;
			3665: Pixel = 193;
			3666: Pixel = 194;
			3667: Pixel = 204;
			3668: Pixel = 206;
			3669: Pixel = 186;
			3670: Pixel = 118;
			3671: Pixel = 80;
			3672: Pixel = 77;
			3673: Pixel = 100;
			3674: Pixel = 124;
			3675: Pixel = 165;
			3676: Pixel = 204;
			3677: Pixel = 88;
			3678: Pixel = 33;
			3679: Pixel = 51;
			3680: Pixel = 49;
			3681: Pixel = 45;
			3682: Pixel = 54;
			3683: Pixel = 50;
			3684: Pixel = 64;
			3685: Pixel = 144;
			3686: Pixel = 146;
			3687: Pixel = 157;
			3688: Pixel = 164;
			3689: Pixel = 160;
			3690: Pixel = 160;
			3691: Pixel = 159;
			3692: Pixel = 158;
			3693: Pixel = 157;
			3694: Pixel = 156;
			3695: Pixel = 155;
			3696: Pixel = 154;
			3697: Pixel = 154;
			3698: Pixel = 153;
			3699: Pixel = 153;
			3700: Pixel = 106;
			3701: Pixel = 103;
			3702: Pixel = 100;
			3703: Pixel = 99;
			3704: Pixel = 106;
			3705: Pixel = 129;
			3706: Pixel = 153;
			3707: Pixel = 168;
			3708: Pixel = 170;
			3709: Pixel = 171;
			3710: Pixel = 168;
			3711: Pixel = 146;
			3712: Pixel = 96;
			3713: Pixel = 73;
			3714: Pixel = 87;
			3715: Pixel = 94;
			3716: Pixel = 97;
			3717: Pixel = 98;
			3718: Pixel = 99;
			3719: Pixel = 98;
			3720: Pixel = 98;
			3721: Pixel = 100;
			3722: Pixel = 87;
			3723: Pixel = 113;
			3724: Pixel = 208;
			3725: Pixel = 195;
			3726: Pixel = 163;
			3727: Pixel = 134;
			3728: Pixel = 148;
			3729: Pixel = 115;
			3730: Pixel = 115;
			3731: Pixel = 137;
			3732: Pixel = 129;
			3733: Pixel = 119;
			3734: Pixel = 128;
			3735: Pixel = 130;
			3736: Pixel = 123;
			3737: Pixel = 135;
			3738: Pixel = 141;
			3739: Pixel = 119;
			3740: Pixel = 126;
			3741: Pixel = 89;
			3742: Pixel = 77;
			3743: Pixel = 73;
			3744: Pixel = 58;
			3745: Pixel = 43;
			3746: Pixel = 95;
			3747: Pixel = 109;
			3748: Pixel = 53;
			3749: Pixel = 82;
			3750: Pixel = 92;
			3751: Pixel = 59;
			3752: Pixel = 63;
			3753: Pixel = 60;
			3754: Pixel = 133;
			3755: Pixel = 154;
			3756: Pixel = 176;
			3757: Pixel = 189;
			3758: Pixel = 179;
			3759: Pixel = 187;
			3760: Pixel = 188;
			3761: Pixel = 186;
			3762: Pixel = 187;
			3763: Pixel = 190;
			3764: Pixel = 191;
			3765: Pixel = 197;
			3766: Pixel = 206;
			3767: Pixel = 178;
			3768: Pixel = 121;
			3769: Pixel = 118;
			3770: Pixel = 122;
			3771: Pixel = 117;
			3772: Pixel = 140;
			3773: Pixel = 157;
			3774: Pixel = 171;
			3775: Pixel = 199;
			3776: Pixel = 95;
			3777: Pixel = 32;
			3778: Pixel = 54;
			3779: Pixel = 54;
			3780: Pixel = 49;
			3781: Pixel = 44;
			3782: Pixel = 56;
			3783: Pixel = 50;
			3784: Pixel = 106;
			3785: Pixel = 151;
			3786: Pixel = 147;
			3787: Pixel = 164;
			3788: Pixel = 163;
			3789: Pixel = 162;
			3790: Pixel = 161;
			3791: Pixel = 160;
			3792: Pixel = 159;
			3793: Pixel = 158;
			3794: Pixel = 156;
			3795: Pixel = 155;
			3796: Pixel = 155;
			3797: Pixel = 155;
			3798: Pixel = 154;
			3799: Pixel = 151;
			3800: Pixel = 106;
			3801: Pixel = 104;
			3802: Pixel = 102;
			3803: Pixel = 100;
			3804: Pixel = 104;
			3805: Pixel = 127;
			3806: Pixel = 153;
			3807: Pixel = 169;
			3808: Pixel = 171;
			3809: Pixel = 171;
			3810: Pixel = 168;
			3811: Pixel = 146;
			3812: Pixel = 98;
			3813: Pixel = 73;
			3814: Pixel = 88;
			3815: Pixel = 94;
			3816: Pixel = 96;
			3817: Pixel = 99;
			3818: Pixel = 99;
			3819: Pixel = 97;
			3820: Pixel = 97;
			3821: Pixel = 101;
			3822: Pixel = 98;
			3823: Pixel = 88;
			3824: Pixel = 194;
			3825: Pixel = 202;
			3826: Pixel = 181;
			3827: Pixel = 159;
			3828: Pixel = 132;
			3829: Pixel = 109;
			3830: Pixel = 135;
			3831: Pixel = 133;
			3832: Pixel = 112;
			3833: Pixel = 123;
			3834: Pixel = 127;
			3835: Pixel = 121;
			3836: Pixel = 131;
			3837: Pixel = 118;
			3838: Pixel = 122;
			3839: Pixel = 117;
			3840: Pixel = 74;
			3841: Pixel = 71;
			3842: Pixel = 68;
			3843: Pixel = 53;
			3844: Pixel = 46;
			3845: Pixel = 60;
			3846: Pixel = 98;
			3847: Pixel = 56;
			3848: Pixel = 82;
			3849: Pixel = 105;
			3850: Pixel = 67;
			3851: Pixel = 44;
			3852: Pixel = 93;
			3853: Pixel = 140;
			3854: Pixel = 149;
			3855: Pixel = 187;
			3856: Pixel = 192;
			3857: Pixel = 177;
			3858: Pixel = 183;
			3859: Pixel = 182;
			3860: Pixel = 178;
			3861: Pixel = 181;
			3862: Pixel = 188;
			3863: Pixel = 191;
			3864: Pixel = 194;
			3865: Pixel = 189;
			3866: Pixel = 122;
			3867: Pixel = 81;
			3868: Pixel = 103;
			3869: Pixel = 114;
			3870: Pixel = 157;
			3871: Pixel = 170;
			3872: Pixel = 168;
			3873: Pixel = 177;
			3874: Pixel = 199;
			3875: Pixel = 102;
			3876: Pixel = 28;
			3877: Pixel = 51;
			3878: Pixel = 54;
			3879: Pixel = 53;
			3880: Pixel = 47;
			3881: Pixel = 50;
			3882: Pixel = 49;
			3883: Pixel = 58;
			3884: Pixel = 137;
			3885: Pixel = 146;
			3886: Pixel = 155;
			3887: Pixel = 166;
			3888: Pixel = 164;
			3889: Pixel = 164;
			3890: Pixel = 162;
			3891: Pixel = 161;
			3892: Pixel = 158;
			3893: Pixel = 158;
			3894: Pixel = 156;
			3895: Pixel = 155;
			3896: Pixel = 155;
			3897: Pixel = 155;
			3898: Pixel = 153;
			3899: Pixel = 152;
			3900: Pixel = 107;
			3901: Pixel = 106;
			3902: Pixel = 102;
			3903: Pixel = 99;
			3904: Pixel = 101;
			3905: Pixel = 123;
			3906: Pixel = 153;
			3907: Pixel = 170;
			3908: Pixel = 171;
			3909: Pixel = 172;
			3910: Pixel = 168;
			3911: Pixel = 148;
			3912: Pixel = 98;
			3913: Pixel = 71;
			3914: Pixel = 87;
			3915: Pixel = 93;
			3916: Pixel = 96;
			3917: Pixel = 97;
			3918: Pixel = 97;
			3919: Pixel = 96;
			3920: Pixel = 97;
			3921: Pixel = 103;
			3922: Pixel = 106;
			3923: Pixel = 86;
			3924: Pixel = 142;
			3925: Pixel = 219;
			3926: Pixel = 174;
			3927: Pixel = 176;
			3928: Pixel = 123;
			3929: Pixel = 125;
			3930: Pixel = 131;
			3931: Pixel = 114;
			3932: Pixel = 126;
			3933: Pixel = 126;
			3934: Pixel = 119;
			3935: Pixel = 129;
			3936: Pixel = 134;
			3937: Pixel = 112;
			3938: Pixel = 76;
			3939: Pixel = 73;
			3940: Pixel = 77;
			3941: Pixel = 68;
			3942: Pixel = 56;
			3943: Pixel = 78;
			3944: Pixel = 37;
			3945: Pixel = 82;
			3946: Pixel = 55;
			3947: Pixel = 52;
			3948: Pixel = 77;
			3949: Pixel = 74;
			3950: Pixel = 82;
			3951: Pixel = 79;
			3952: Pixel = 126;
			3953: Pixel = 149;
			3954: Pixel = 192;
			3955: Pixel = 195;
			3956: Pixel = 183;
			3957: Pixel = 179;
			3958: Pixel = 182;
			3959: Pixel = 175;
			3960: Pixel = 175;
			3961: Pixel = 180;
			3962: Pixel = 189;
			3963: Pixel = 188;
			3964: Pixel = 192;
			3965: Pixel = 119;
			3966: Pixel = 60;
			3967: Pixel = 95;
			3968: Pixel = 118;
			3969: Pixel = 119;
			3970: Pixel = 134;
			3971: Pixel = 163;
			3972: Pixel = 185;
			3973: Pixel = 182;
			3974: Pixel = 85;
			3975: Pixel = 32;
			3976: Pixel = 48;
			3977: Pixel = 51;
			3978: Pixel = 56;
			3979: Pixel = 53;
			3980: Pixel = 46;
			3981: Pixel = 50;
			3982: Pixel = 48;
			3983: Pixel = 89;
			3984: Pixel = 140;
			3985: Pixel = 142;
			3986: Pixel = 165;
			3987: Pixel = 166;
			3988: Pixel = 164;
			3989: Pixel = 163;
			3990: Pixel = 163;
			3991: Pixel = 162;
			3992: Pixel = 160;
			3993: Pixel = 158;
			3994: Pixel = 157;
			3995: Pixel = 157;
			3996: Pixel = 156;
			3997: Pixel = 155;
			3998: Pixel = 153;
			3999: Pixel = 152;
			4000: Pixel = 108;
			4001: Pixel = 106;
			4002: Pixel = 103;
			4003: Pixel = 99;
			4004: Pixel = 96;
			4005: Pixel = 119;
			4006: Pixel = 153;
			4007: Pixel = 169;
			4008: Pixel = 172;
			4009: Pixel = 174;
			4010: Pixel = 169;
			4011: Pixel = 147;
			4012: Pixel = 97;
			4013: Pixel = 71;
			4014: Pixel = 84;
			4015: Pixel = 92;
			4016: Pixel = 97;
			4017: Pixel = 96;
			4018: Pixel = 98;
			4019: Pixel = 98;
			4020: Pixel = 99;
			4021: Pixel = 104;
			4022: Pixel = 108;
			4023: Pixel = 103;
			4024: Pixel = 88;
			4025: Pixel = 186;
			4026: Pixel = 201;
			4027: Pixel = 174;
			4028: Pixel = 130;
			4029: Pixel = 126;
			4030: Pixel = 119;
			4031: Pixel = 122;
			4032: Pixel = 130;
			4033: Pixel = 123;
			4034: Pixel = 124;
			4035: Pixel = 126;
			4036: Pixel = 115;
			4037: Pixel = 90;
			4038: Pixel = 82;
			4039: Pixel = 85;
			4040: Pixel = 77;
			4041: Pixel = 36;
			4042: Pixel = 73;
			4043: Pixel = 75;
			4044: Pixel = 48;
			4045: Pixel = 68;
			4046: Pixel = 57;
			4047: Pixel = 65;
			4048: Pixel = 66;
			4049: Pixel = 71;
			4050: Pixel = 102;
			4051: Pixel = 121;
			4052: Pixel = 128;
			4053: Pixel = 190;
			4054: Pixel = 193;
			4055: Pixel = 186;
			4056: Pixel = 179;
			4057: Pixel = 178;
			4058: Pixel = 178;
			4059: Pixel = 172;
			4060: Pixel = 180;
			4061: Pixel = 182;
			4062: Pixel = 184;
			4063: Pixel = 186;
			4064: Pixel = 197;
			4065: Pixel = 157;
			4066: Pixel = 89;
			4067: Pixel = 99;
			4068: Pixel = 103;
			4069: Pixel = 124;
			4070: Pixel = 130;
			4071: Pixel = 175;
			4072: Pixel = 155;
			4073: Pixel = 61;
			4074: Pixel = 34;
			4075: Pixel = 48;
			4076: Pixel = 54;
			4077: Pixel = 52;
			4078: Pixel = 56;
			4079: Pixel = 47;
			4080: Pixel = 47;
			4081: Pixel = 51;
			4082: Pixel = 58;
			4083: Pixel = 116;
			4084: Pixel = 129;
			4085: Pixel = 148;
			4086: Pixel = 170;
			4087: Pixel = 164;
			4088: Pixel = 162;
			4089: Pixel = 163;
			4090: Pixel = 163;
			4091: Pixel = 162;
			4092: Pixel = 161;
			4093: Pixel = 159;
			4094: Pixel = 159;
			4095: Pixel = 158;
			4096: Pixel = 157;
			4097: Pixel = 155;
			4098: Pixel = 153;
			4099: Pixel = 151;
			4100: Pixel = 108;
			4101: Pixel = 105;
			4102: Pixel = 102;
			4103: Pixel = 99;
			4104: Pixel = 92;
			4105: Pixel = 116;
			4106: Pixel = 151;
			4107: Pixel = 169;
			4108: Pixel = 172;
			4109: Pixel = 174;
			4110: Pixel = 171;
			4111: Pixel = 148;
			4112: Pixel = 98;
			4113: Pixel = 69;
			4114: Pixel = 84;
			4115: Pixel = 92;
			4116: Pixel = 97;
			4117: Pixel = 97;
			4118: Pixel = 96;
			4119: Pixel = 97;
			4120: Pixel = 100;
			4121: Pixel = 105;
			4122: Pixel = 111;
			4123: Pixel = 112;
			4124: Pixel = 87;
			4125: Pixel = 149;
			4126: Pixel = 218;
			4127: Pixel = 185;
			4128: Pixel = 133;
			4129: Pixel = 116;
			4130: Pixel = 112;
			4131: Pixel = 126;
			4132: Pixel = 117;
			4133: Pixel = 125;
			4134: Pixel = 124;
			4135: Pixel = 123;
			4136: Pixel = 97;
			4137: Pixel = 63;
			4138: Pixel = 63;
			4139: Pixel = 86;
			4140: Pixel = 69;
			4141: Pixel = 51;
			4142: Pixel = 66;
			4143: Pixel = 84;
			4144: Pixel = 58;
			4145: Pixel = 42;
			4146: Pixel = 52;
			4147: Pixel = 57;
			4148: Pixel = 52;
			4149: Pixel = 83;
			4150: Pixel = 86;
			4151: Pixel = 125;
			4152: Pixel = 166;
			4153: Pixel = 179;
			4154: Pixel = 181;
			4155: Pixel = 175;
			4156: Pixel = 171;
			4157: Pixel = 175;
			4158: Pixel = 175;
			4159: Pixel = 173;
			4160: Pixel = 175;
			4161: Pixel = 191;
			4162: Pixel = 193;
			4163: Pixel = 195;
			4164: Pixel = 199;
			4165: Pixel = 189;
			4166: Pixel = 115;
			4167: Pixel = 72;
			4168: Pixel = 82;
			4169: Pixel = 101;
			4170: Pixel = 142;
			4171: Pixel = 149;
			4172: Pixel = 64;
			4173: Pixel = 33;
			4174: Pixel = 48;
			4175: Pixel = 52;
			4176: Pixel = 56;
			4177: Pixel = 57;
			4178: Pixel = 54;
			4179: Pixel = 43;
			4180: Pixel = 50;
			4181: Pixel = 49;
			4182: Pixel = 79;
			4183: Pixel = 131;
			4184: Pixel = 126;
			4185: Pixel = 159;
			4186: Pixel = 168;
			4187: Pixel = 164;
			4188: Pixel = 163;
			4189: Pixel = 163;
			4190: Pixel = 163;
			4191: Pixel = 162;
			4192: Pixel = 161;
			4193: Pixel = 160;
			4194: Pixel = 161;
			4195: Pixel = 158;
			4196: Pixel = 157;
			4197: Pixel = 156;
			4198: Pixel = 154;
			4199: Pixel = 151;
			4200: Pixel = 105;
			4201: Pixel = 105;
			4202: Pixel = 103;
			4203: Pixel = 98;
			4204: Pixel = 90;
			4205: Pixel = 115;
			4206: Pixel = 150;
			4207: Pixel = 168;
			4208: Pixel = 172;
			4209: Pixel = 174;
			4210: Pixel = 170;
			4211: Pixel = 149;
			4212: Pixel = 99;
			4213: Pixel = 71;
			4214: Pixel = 86;
			4215: Pixel = 94;
			4216: Pixel = 98;
			4217: Pixel = 100;
			4218: Pixel = 98;
			4219: Pixel = 98;
			4220: Pixel = 100;
			4221: Pixel = 105;
			4222: Pixel = 112;
			4223: Pixel = 114;
			4224: Pixel = 92;
			4225: Pixel = 146;
			4226: Pixel = 229;
			4227: Pixel = 167;
			4228: Pixel = 109;
			4229: Pixel = 122;
			4230: Pixel = 119;
			4231: Pixel = 113;
			4232: Pixel = 133;
			4233: Pixel = 137;
			4234: Pixel = 115;
			4235: Pixel = 69;
			4236: Pixel = 72;
			4237: Pixel = 61;
			4238: Pixel = 41;
			4239: Pixel = 65;
			4240: Pixel = 79;
			4241: Pixel = 68;
			4242: Pixel = 52;
			4243: Pixel = 91;
			4244: Pixel = 85;
			4245: Pixel = 48;
			4246: Pixel = 47;
			4247: Pixel = 31;
			4248: Pixel = 71;
			4249: Pixel = 104;
			4250: Pixel = 120;
			4251: Pixel = 163;
			4252: Pixel = 181;
			4253: Pixel = 186;
			4254: Pixel = 180;
			4255: Pixel = 161;
			4256: Pixel = 170;
			4257: Pixel = 178;
			4258: Pixel = 164;
			4259: Pixel = 173;
			4260: Pixel = 189;
			4261: Pixel = 199;
			4262: Pixel = 198;
			4263: Pixel = 197;
			4264: Pixel = 200;
			4265: Pixel = 194;
			4266: Pixel = 137;
			4267: Pixel = 66;
			4268: Pixel = 53;
			4269: Pixel = 84;
			4270: Pixel = 136;
			4271: Pixel = 143;
			4272: Pixel = 60;
			4273: Pixel = 43;
			4274: Pixel = 46;
			4275: Pixel = 55;
			4276: Pixel = 57;
			4277: Pixel = 61;
			4278: Pixel = 51;
			4279: Pixel = 44;
			4280: Pixel = 49;
			4281: Pixel = 48;
			4282: Pixel = 110;
			4283: Pixel = 134;
			4284: Pixel = 136;
			4285: Pixel = 159;
			4286: Pixel = 164;
			4287: Pixel = 166;
			4288: Pixel = 165;
			4289: Pixel = 161;
			4290: Pixel = 161;
			4291: Pixel = 162;
			4292: Pixel = 162;
			4293: Pixel = 161;
			4294: Pixel = 160;
			4295: Pixel = 158;
			4296: Pixel = 158;
			4297: Pixel = 157;
			4298: Pixel = 154;
			4299: Pixel = 151;
			4300: Pixel = 103;
			4301: Pixel = 104;
			4302: Pixel = 102;
			4303: Pixel = 99;
			4304: Pixel = 91;
			4305: Pixel = 115;
			4306: Pixel = 150;
			4307: Pixel = 168;
			4308: Pixel = 172;
			4309: Pixel = 174;
			4310: Pixel = 170;
			4311: Pixel = 150;
			4312: Pixel = 101;
			4313: Pixel = 72;
			4314: Pixel = 85;
			4315: Pixel = 94;
			4316: Pixel = 98;
			4317: Pixel = 101;
			4318: Pixel = 100;
			4319: Pixel = 100;
			4320: Pixel = 102;
			4321: Pixel = 107;
			4322: Pixel = 115;
			4323: Pixel = 116;
			4324: Pixel = 100;
			4325: Pixel = 130;
			4326: Pixel = 224;
			4327: Pixel = 130;
			4328: Pixel = 103;
			4329: Pixel = 113;
			4330: Pixel = 117;
			4331: Pixel = 126;
			4332: Pixel = 112;
			4333: Pixel = 107;
			4334: Pixel = 97;
			4335: Pixel = 52;
			4336: Pixel = 68;
			4337: Pixel = 43;
			4338: Pixel = 49;
			4339: Pixel = 52;
			4340: Pixel = 72;
			4341: Pixel = 68;
			4342: Pixel = 64;
			4343: Pixel = 59;
			4344: Pixel = 102;
			4345: Pixel = 58;
			4346: Pixel = 28;
			4347: Pixel = 69;
			4348: Pixel = 130;
			4349: Pixel = 148;
			4350: Pixel = 158;
			4351: Pixel = 156;
			4352: Pixel = 183;
			4353: Pixel = 186;
			4354: Pixel = 169;
			4355: Pixel = 162;
			4356: Pixel = 174;
			4357: Pixel = 165;
			4358: Pixel = 167;
			4359: Pixel = 185;
			4360: Pixel = 195;
			4361: Pixel = 198;
			4362: Pixel = 200;
			4363: Pixel = 202;
			4364: Pixel = 208;
			4365: Pixel = 206;
			4366: Pixel = 157;
			4367: Pixel = 80;
			4368: Pixel = 41;
			4369: Pixel = 62;
			4370: Pixel = 133;
			4371: Pixel = 146;
			4372: Pixel = 47;
			4373: Pixel = 47;
			4374: Pixel = 51;
			4375: Pixel = 54;
			4376: Pixel = 59;
			4377: Pixel = 60;
			4378: Pixel = 46;
			4379: Pixel = 48;
			4380: Pixel = 46;
			4381: Pixel = 66;
			4382: Pixel = 134;
			4383: Pixel = 134;
			4384: Pixel = 151;
			4385: Pixel = 151;
			4386: Pixel = 153;
			4387: Pixel = 159;
			4388: Pixel = 162;
			4389: Pixel = 161;
			4390: Pixel = 161;
			4391: Pixel = 161;
			4392: Pixel = 163;
			4393: Pixel = 161;
			4394: Pixel = 159;
			4395: Pixel = 157;
			4396: Pixel = 157;
			4397: Pixel = 157;
			4398: Pixel = 155;
			4399: Pixel = 151;
			4400: Pixel = 104;
			4401: Pixel = 103;
			4402: Pixel = 101;
			4403: Pixel = 99;
			4404: Pixel = 92;
			4405: Pixel = 114;
			4406: Pixel = 150;
			4407: Pixel = 168;
			4408: Pixel = 173;
			4409: Pixel = 174;
			4410: Pixel = 172;
			4411: Pixel = 149;
			4412: Pixel = 103;
			4413: Pixel = 74;
			4414: Pixel = 85;
			4415: Pixel = 96;
			4416: Pixel = 101;
			4417: Pixel = 103;
			4418: Pixel = 102;
			4419: Pixel = 100;
			4420: Pixel = 98;
			4421: Pixel = 122;
			4422: Pixel = 121;
			4423: Pixel = 114;
			4424: Pixel = 112;
			4425: Pixel = 108;
			4426: Pixel = 198;
			4427: Pixel = 131;
			4428: Pixel = 112;
			4429: Pixel = 111;
			4430: Pixel = 125;
			4431: Pixel = 130;
			4432: Pixel = 103;
			4433: Pixel = 70;
			4434: Pixel = 51;
			4435: Pixel = 61;
			4436: Pixel = 67;
			4437: Pixel = 48;
			4438: Pixel = 58;
			4439: Pixel = 49;
			4440: Pixel = 53;
			4441: Pixel = 55;
			4442: Pixel = 87;
			4443: Pixel = 79;
			4444: Pixel = 89;
			4445: Pixel = 31;
			4446: Pixel = 56;
			4447: Pixel = 133;
			4448: Pixel = 152;
			4449: Pixel = 180;
			4450: Pixel = 160;
			4451: Pixel = 155;
			4452: Pixel = 182;
			4453: Pixel = 183;
			4454: Pixel = 168;
			4455: Pixel = 167;
			4456: Pixel = 156;
			4457: Pixel = 162;
			4458: Pixel = 178;
			4459: Pixel = 190;
			4460: Pixel = 196;
			4461: Pixel = 200;
			4462: Pixel = 201;
			4463: Pixel = 206;
			4464: Pixel = 210;
			4465: Pixel = 211;
			4466: Pixel = 178;
			4467: Pixel = 97;
			4468: Pixel = 43;
			4469: Pixel = 41;
			4470: Pixel = 108;
			4471: Pixel = 155;
			4472: Pixel = 58;
			4473: Pixel = 50;
			4474: Pixel = 55;
			4475: Pixel = 57;
			4476: Pixel = 63;
			4477: Pixel = 56;
			4478: Pixel = 44;
			4479: Pixel = 54;
			4480: Pixel = 42;
			4481: Pixel = 91;
			4482: Pixel = 142;
			4483: Pixel = 141;
			4484: Pixel = 162;
			4485: Pixel = 153;
			4486: Pixel = 150;
			4487: Pixel = 149;
			4488: Pixel = 149;
			4489: Pixel = 152;
			4490: Pixel = 155;
			4491: Pixel = 157;
			4492: Pixel = 160;
			4493: Pixel = 161;
			4494: Pixel = 160;
			4495: Pixel = 158;
			4496: Pixel = 156;
			4497: Pixel = 155;
			4498: Pixel = 154;
			4499: Pixel = 151;
			4500: Pixel = 105;
			4501: Pixel = 102;
			4502: Pixel = 99;
			4503: Pixel = 96;
			4504: Pixel = 90;
			4505: Pixel = 113;
			4506: Pixel = 148;
			4507: Pixel = 168;
			4508: Pixel = 174;
			4509: Pixel = 174;
			4510: Pixel = 171;
			4511: Pixel = 149;
			4512: Pixel = 102;
			4513: Pixel = 77;
			4514: Pixel = 91;
			4515: Pixel = 97;
			4516: Pixel = 100;
			4517: Pixel = 102;
			4518: Pixel = 102;
			4519: Pixel = 101;
			4520: Pixel = 103;
			4521: Pixel = 115;
			4522: Pixel = 114;
			4523: Pixel = 118;
			4524: Pixel = 121;
			4525: Pixel = 107;
			4526: Pixel = 156;
			4527: Pixel = 146;
			4528: Pixel = 109;
			4529: Pixel = 130;
			4530: Pixel = 131;
			4531: Pixel = 118;
			4532: Pixel = 73;
			4533: Pixel = 65;
			4534: Pixel = 53;
			4535: Pixel = 43;
			4536: Pixel = 70;
			4537: Pixel = 54;
			4538: Pixel = 58;
			4539: Pixel = 49;
			4540: Pixel = 59;
			4541: Pixel = 51;
			4542: Pixel = 74;
			4543: Pixel = 67;
			4544: Pixel = 86;
			4545: Pixel = 69;
			4546: Pixel = 120;
			4547: Pixel = 145;
			4548: Pixel = 175;
			4549: Pixel = 186;
			4550: Pixel = 171;
			4551: Pixel = 149;
			4552: Pixel = 190;
			4553: Pixel = 174;
			4554: Pixel = 159;
			4555: Pixel = 155;
			4556: Pixel = 162;
			4557: Pixel = 171;
			4558: Pixel = 179;
			4559: Pixel = 192;
			4560: Pixel = 196;
			4561: Pixel = 201;
			4562: Pixel = 203;
			4563: Pixel = 206;
			4564: Pixel = 210;
			4565: Pixel = 214;
			4566: Pixel = 193;
			4567: Pixel = 114;
			4568: Pixel = 54;
			4569: Pixel = 36;
			4570: Pixel = 88;
			4571: Pixel = 156;
			4572: Pixel = 65;
			4573: Pixel = 48;
			4574: Pixel = 57;
			4575: Pixel = 58;
			4576: Pixel = 61;
			4577: Pixel = 53;
			4578: Pixel = 48;
			4579: Pixel = 51;
			4580: Pixel = 49;
			4581: Pixel = 126;
			4582: Pixel = 139;
			4583: Pixel = 153;
			4584: Pixel = 165;
			4585: Pixel = 161;
			4586: Pixel = 157;
			4587: Pixel = 154;
			4588: Pixel = 151;
			4589: Pixel = 150;
			4590: Pixel = 147;
			4591: Pixel = 145;
			4592: Pixel = 148;
			4593: Pixel = 152;
			4594: Pixel = 154;
			4595: Pixel = 154;
			4596: Pixel = 154;
			4597: Pixel = 153;
			4598: Pixel = 153;
			4599: Pixel = 150;
			4600: Pixel = 102;
			4601: Pixel = 102;
			4602: Pixel = 99;
			4603: Pixel = 97;
			4604: Pixel = 89;
			4605: Pixel = 113;
			4606: Pixel = 150;
			4607: Pixel = 169;
			4608: Pixel = 174;
			4609: Pixel = 175;
			4610: Pixel = 171;
			4611: Pixel = 150;
			4612: Pixel = 100;
			4613: Pixel = 75;
			4614: Pixel = 89;
			4615: Pixel = 97;
			4616: Pixel = 100;
			4617: Pixel = 102;
			4618: Pixel = 104;
			4619: Pixel = 102;
			4620: Pixel = 105;
			4621: Pixel = 112;
			4622: Pixel = 117;
			4623: Pixel = 117;
			4624: Pixel = 111;
			4625: Pixel = 117;
			4626: Pixel = 124;
			4627: Pixel = 125;
			4628: Pixel = 123;
			4629: Pixel = 133;
			4630: Pixel = 127;
			4631: Pixel = 79;
			4632: Pixel = 50;
			4633: Pixel = 61;
			4634: Pixel = 67;
			4635: Pixel = 44;
			4636: Pixel = 59;
			4637: Pixel = 80;
			4638: Pixel = 52;
			4639: Pixel = 46;
			4640: Pixel = 63;
			4641: Pixel = 58;
			4642: Pixel = 60;
			4643: Pixel = 59;
			4644: Pixel = 37;
			4645: Pixel = 118;
			4646: Pixel = 138;
			4647: Pixel = 163;
			4648: Pixel = 164;
			4649: Pixel = 187;
			4650: Pixel = 177;
			4651: Pixel = 166;
			4652: Pixel = 183;
			4653: Pixel = 159;
			4654: Pixel = 160;
			4655: Pixel = 161;
			4656: Pixel = 170;
			4657: Pixel = 174;
			4658: Pixel = 178;
			4659: Pixel = 188;
			4660: Pixel = 196;
			4661: Pixel = 197;
			4662: Pixel = 200;
			4663: Pixel = 204;
			4664: Pixel = 208;
			4665: Pixel = 212;
			4666: Pixel = 203;
			4667: Pixel = 137;
			4668: Pixel = 71;
			4669: Pixel = 36;
			4670: Pixel = 70;
			4671: Pixel = 154;
			4672: Pixel = 74;
			4673: Pixel = 48;
			4674: Pixel = 59;
			4675: Pixel = 61;
			4676: Pixel = 60;
			4677: Pixel = 49;
			4678: Pixel = 53;
			4679: Pixel = 44;
			4680: Pixel = 77;
			4681: Pixel = 140;
			4682: Pixel = 137;
			4683: Pixel = 161;
			4684: Pixel = 163;
			4685: Pixel = 160;
			4686: Pixel = 161;
			4687: Pixel = 163;
			4688: Pixel = 162;
			4689: Pixel = 158;
			4690: Pixel = 154;
			4691: Pixel = 146;
			4692: Pixel = 146;
			4693: Pixel = 144;
			4694: Pixel = 143;
			4695: Pixel = 144;
			4696: Pixel = 147;
			4697: Pixel = 151;
			4698: Pixel = 153;
			4699: Pixel = 151;
			4700: Pixel = 101;
			4701: Pixel = 100;
			4702: Pixel = 98;
			4703: Pixel = 97;
			4704: Pixel = 90;
			4705: Pixel = 112;
			4706: Pixel = 150;
			4707: Pixel = 168;
			4708: Pixel = 173;
			4709: Pixel = 176;
			4710: Pixel = 171;
			4711: Pixel = 149;
			4712: Pixel = 101;
			4713: Pixel = 75;
			4714: Pixel = 87;
			4715: Pixel = 97;
			4716: Pixel = 101;
			4717: Pixel = 102;
			4718: Pixel = 102;
			4719: Pixel = 102;
			4720: Pixel = 105;
			4721: Pixel = 112;
			4722: Pixel = 118;
			4723: Pixel = 117;
			4724: Pixel = 125;
			4725: Pixel = 143;
			4726: Pixel = 101;
			4727: Pixel = 121;
			4728: Pixel = 130;
			4729: Pixel = 127;
			4730: Pixel = 104;
			4731: Pixel = 71;
			4732: Pixel = 61;
			4733: Pixel = 66;
			4734: Pixel = 67;
			4735: Pixel = 44;
			4736: Pixel = 74;
			4737: Pixel = 64;
			4738: Pixel = 41;
			4739: Pixel = 55;
			4740: Pixel = 54;
			4741: Pixel = 67;
			4742: Pixel = 69;
			4743: Pixel = 47;
			4744: Pixel = 85;
			4745: Pixel = 125;
			4746: Pixel = 168;
			4747: Pixel = 172;
			4748: Pixel = 159;
			4749: Pixel = 184;
			4750: Pixel = 194;
			4751: Pixel = 162;
			4752: Pixel = 118;
			4753: Pixel = 135;
			4754: Pixel = 154;
			4755: Pixel = 170;
			4756: Pixel = 181;
			4757: Pixel = 179;
			4758: Pixel = 176;
			4759: Pixel = 181;
			4760: Pixel = 192;
			4761: Pixel = 194;
			4762: Pixel = 195;
			4763: Pixel = 200;
			4764: Pixel = 205;
			4765: Pixel = 214;
			4766: Pixel = 210;
			4767: Pixel = 140;
			4768: Pixel = 58;
			4769: Pixel = 38;
			4770: Pixel = 55;
			4771: Pixel = 150;
			4772: Pixel = 91;
			4773: Pixel = 56;
			4774: Pixel = 60;
			4775: Pixel = 65;
			4776: Pixel = 57;
			4777: Pixel = 49;
			4778: Pixel = 53;
			4779: Pixel = 45;
			4780: Pixel = 108;
			4781: Pixel = 137;
			4782: Pixel = 142;
			4783: Pixel = 163;
			4784: Pixel = 161;
			4785: Pixel = 160;
			4786: Pixel = 159;
			4787: Pixel = 162;
			4788: Pixel = 165;
			4789: Pixel = 162;
			4790: Pixel = 157;
			4791: Pixel = 154;
			4792: Pixel = 150;
			4793: Pixel = 146;
			4794: Pixel = 144;
			4795: Pixel = 143;
			4796: Pixel = 141;
			4797: Pixel = 142;
			4798: Pixel = 144;
			4799: Pixel = 145;
			4800: Pixel = 101;
			4801: Pixel = 100;
			4802: Pixel = 100;
			4803: Pixel = 100;
			4804: Pixel = 91;
			4805: Pixel = 111;
			4806: Pixel = 150;
			4807: Pixel = 168;
			4808: Pixel = 175;
			4809: Pixel = 176;
			4810: Pixel = 172;
			4811: Pixel = 151;
			4812: Pixel = 101;
			4813: Pixel = 76;
			4814: Pixel = 88;
			4815: Pixel = 95;
			4816: Pixel = 102;
			4817: Pixel = 102;
			4818: Pixel = 101;
			4819: Pixel = 102;
			4820: Pixel = 104;
			4821: Pixel = 113;
			4822: Pixel = 118;
			4823: Pixel = 115;
			4824: Pixel = 154;
			4825: Pixel = 121;
			4826: Pixel = 19;
			4827: Pixel = 82;
			4828: Pixel = 159;
			4829: Pixel = 99;
			4830: Pixel = 65;
			4831: Pixel = 82;
			4832: Pixel = 49;
			4833: Pixel = 96;
			4834: Pixel = 56;
			4835: Pixel = 47;
			4836: Pixel = 61;
			4837: Pixel = 53;
			4838: Pixel = 46;
			4839: Pixel = 50;
			4840: Pixel = 71;
			4841: Pixel = 75;
			4842: Pixel = 50;
			4843: Pixel = 66;
			4844: Pixel = 128;
			4845: Pixel = 160;
			4846: Pixel = 185;
			4847: Pixel = 175;
			4848: Pixel = 159;
			4849: Pixel = 198;
			4850: Pixel = 170;
			4851: Pixel = 126;
			4852: Pixel = 126;
			4853: Pixel = 117;
			4854: Pixel = 90;
			4855: Pixel = 97;
			4856: Pixel = 140;
			4857: Pixel = 176;
			4858: Pixel = 175;
			4859: Pixel = 175;
			4860: Pixel = 188;
			4861: Pixel = 192;
			4862: Pixel = 189;
			4863: Pixel = 196;
			4864: Pixel = 199;
			4865: Pixel = 180;
			4866: Pixel = 140;
			4867: Pixel = 99;
			4868: Pixel = 57;
			4869: Pixel = 40;
			4870: Pixel = 46;
			4871: Pixel = 140;
			4872: Pixel = 109;
			4873: Pixel = 51;
			4874: Pixel = 65;
			4875: Pixel = 64;
			4876: Pixel = 52;
			4877: Pixel = 50;
			4878: Pixel = 52;
			4879: Pixel = 56;
			4880: Pixel = 128;
			4881: Pixel = 134;
			4882: Pixel = 153;
			4883: Pixel = 162;
			4884: Pixel = 157;
			4885: Pixel = 158;
			4886: Pixel = 157;
			4887: Pixel = 156;
			4888: Pixel = 159;
			4889: Pixel = 160;
			4890: Pixel = 155;
			4891: Pixel = 154;
			4892: Pixel = 154;
			4893: Pixel = 153;
			4894: Pixel = 153;
			4895: Pixel = 150;
			4896: Pixel = 143;
			4897: Pixel = 141;
			4898: Pixel = 138;
			4899: Pixel = 133;
			4900: Pixel = 101;
			4901: Pixel = 103;
			4902: Pixel = 103;
			4903: Pixel = 99;
			4904: Pixel = 88;
			4905: Pixel = 110;
			4906: Pixel = 148;
			4907: Pixel = 169;
			4908: Pixel = 174;
			4909: Pixel = 176;
			4910: Pixel = 174;
			4911: Pixel = 152;
			4912: Pixel = 102;
			4913: Pixel = 76;
			4914: Pixel = 89;
			4915: Pixel = 98;
			4916: Pixel = 103;
			4917: Pixel = 101;
			4918: Pixel = 99;
			4919: Pixel = 100;
			4920: Pixel = 103;
			4921: Pixel = 103;
			4922: Pixel = 111;
			4923: Pixel = 143;
			4924: Pixel = 150;
			4925: Pixel = 134;
			4926: Pixel = 88;
			4927: Pixel = 107;
			4928: Pixel = 109;
			4929: Pixel = 59;
			4930: Pixel = 75;
			4931: Pixel = 77;
			4932: Pixel = 69;
			4933: Pixel = 76;
			4934: Pixel = 65;
			4935: Pixel = 54;
			4936: Pixel = 52;
			4937: Pixel = 79;
			4938: Pixel = 46;
			4939: Pixel = 34;
			4940: Pixel = 62;
			4941: Pixel = 68;
			4942: Pixel = 41;
			4943: Pixel = 117;
			4944: Pixel = 159;
			4945: Pixel = 177;
			4946: Pixel = 193;
			4947: Pixel = 167;
			4948: Pixel = 188;
			4949: Pixel = 153;
			4950: Pixel = 113;
			4951: Pixel = 130;
			4952: Pixel = 123;
			4953: Pixel = 137;
			4954: Pixel = 109;
			4955: Pixel = 93;
			4956: Pixel = 83;
			4957: Pixel = 129;
			4958: Pixel = 164;
			4959: Pixel = 167;
			4960: Pixel = 185;
			4961: Pixel = 192;
			4962: Pixel = 189;
			4963: Pixel = 185;
			4964: Pixel = 139;
			4965: Pixel = 97;
			4966: Pixel = 91;
			4967: Pixel = 104;
			4968: Pixel = 82;
			4969: Pixel = 49;
			4970: Pixel = 41;
			4971: Pixel = 130;
			4972: Pixel = 122;
			4973: Pixel = 49;
			4974: Pixel = 67;
			4975: Pixel = 60;
			4976: Pixel = 49;
			4977: Pixel = 53;
			4978: Pixel = 50;
			4979: Pixel = 78;
			4980: Pixel = 136;
			4981: Pixel = 135;
			4982: Pixel = 160;
			4983: Pixel = 159;
			4984: Pixel = 157;
			4985: Pixel = 156;
			4986: Pixel = 155;
			4987: Pixel = 154;
			4988: Pixel = 156;
			4989: Pixel = 157;
			4990: Pixel = 155;
			4991: Pixel = 153;
			4992: Pixel = 153;
			4993: Pixel = 155;
			4994: Pixel = 157;
			4995: Pixel = 154;
			4996: Pixel = 149;
			4997: Pixel = 147;
			4998: Pixel = 139;
			4999: Pixel = 133;
			5000: Pixel = 100;
			5001: Pixel = 100;
			5002: Pixel = 99;
			5003: Pixel = 96;
			5004: Pixel = 84;
			5005: Pixel = 108;
			5006: Pixel = 148;
			5007: Pixel = 169;
			5008: Pixel = 176;
			5009: Pixel = 177;
			5010: Pixel = 172;
			5011: Pixel = 153;
			5012: Pixel = 105;
			5013: Pixel = 74;
			5014: Pixel = 85;
			5015: Pixel = 95;
			5016: Pixel = 101;
			5017: Pixel = 100;
			5018: Pixel = 98;
			5019: Pixel = 97;
			5020: Pixel = 94;
			5021: Pixel = 129;
			5022: Pixel = 149;
			5023: Pixel = 149;
			5024: Pixel = 156;
			5025: Pixel = 149;
			5026: Pixel = 134;
			5027: Pixel = 70;
			5028: Pixel = 55;
			5029: Pixel = 77;
			5030: Pixel = 100;
			5031: Pixel = 77;
			5032: Pixel = 94;
			5033: Pixel = 48;
			5034: Pixel = 66;
			5035: Pixel = 66;
			5036: Pixel = 40;
			5037: Pixel = 59;
			5038: Pixel = 85;
			5039: Pixel = 46;
			5040: Pixel = 41;
			5041: Pixel = 31;
			5042: Pixel = 87;
			5043: Pixel = 149;
			5044: Pixel = 174;
			5045: Pixel = 187;
			5046: Pixel = 195;
			5047: Pixel = 189;
			5048: Pixel = 127;
			5049: Pixel = 65;
			5050: Pixel = 65;
			5051: Pixel = 55;
			5052: Pixel = 50;
			5053: Pixel = 58;
			5054: Pixel = 43;
			5055: Pixel = 95;
			5056: Pixel = 131;
			5057: Pixel = 125;
			5058: Pixel = 146;
			5059: Pixel = 159;
			5060: Pixel = 184;
			5061: Pixel = 198;
			5062: Pixel = 198;
			5063: Pixel = 131;
			5064: Pixel = 74;
			5065: Pixel = 60;
			5066: Pixel = 52;
			5067: Pixel = 60;
			5068: Pixel = 64;
			5069: Pixel = 48;
			5070: Pixel = 41;
			5071: Pixel = 124;
			5072: Pixel = 130;
			5073: Pixel = 56;
			5074: Pixel = 65;
			5075: Pixel = 54;
			5076: Pixel = 47;
			5077: Pixel = 54;
			5078: Pixel = 41;
			5079: Pixel = 101;
			5080: Pixel = 140;
			5081: Pixel = 144;
			5082: Pixel = 161;
			5083: Pixel = 156;
			5084: Pixel = 154;
			5085: Pixel = 155;
			5086: Pixel = 155;
			5087: Pixel = 155;
			5088: Pixel = 155;
			5089: Pixel = 156;
			5090: Pixel = 154;
			5091: Pixel = 153;
			5092: Pixel = 153;
			5093: Pixel = 153;
			5094: Pixel = 154;
			5095: Pixel = 152;
			5096: Pixel = 146;
			5097: Pixel = 146;
			5098: Pixel = 142;
			5099: Pixel = 137;
			5100: Pixel = 97;
			5101: Pixel = 95;
			5102: Pixel = 93;
			5103: Pixel = 90;
			5104: Pixel = 77;
			5105: Pixel = 101;
			5106: Pixel = 147;
			5107: Pixel = 170;
			5108: Pixel = 176;
			5109: Pixel = 177;
			5110: Pixel = 172;
			5111: Pixel = 150;
			5112: Pixel = 103;
			5113: Pixel = 72;
			5114: Pixel = 87;
			5115: Pixel = 94;
			5116: Pixel = 98;
			5117: Pixel = 97;
			5118: Pixel = 96;
			5119: Pixel = 89;
			5120: Pixel = 105;
			5121: Pixel = 195;
			5122: Pixel = 147;
			5123: Pixel = 140;
			5124: Pixel = 151;
			5125: Pixel = 118;
			5126: Pixel = 50;
			5127: Pixel = 46;
			5128: Pixel = 79;
			5129: Pixel = 79;
			5130: Pixel = 63;
			5131: Pixel = 92;
			5132: Pixel = 96;
			5133: Pixel = 47;
			5134: Pixel = 48;
			5135: Pixel = 75;
			5136: Pixel = 59;
			5137: Pixel = 35;
			5138: Pixel = 72;
			5139: Pixel = 72;
			5140: Pixel = 42;
			5141: Pixel = 53;
			5142: Pixel = 131;
			5143: Pixel = 172;
			5144: Pixel = 176;
			5145: Pixel = 195;
			5146: Pixel = 202;
			5147: Pixel = 129;
			5148: Pixel = 52;
			5149: Pixel = 49;
			5150: Pixel = 56;
			5151: Pixel = 46;
			5152: Pixel = 60;
			5153: Pixel = 152;
			5154: Pixel = 95;
			5155: Pixel = 49;
			5156: Pixel = 116;
			5157: Pixel = 130;
			5158: Pixel = 138;
			5159: Pixel = 153;
			5160: Pixel = 186;
			5161: Pixel = 218;
			5162: Pixel = 132;
			5163: Pixel = 40;
			5164: Pixel = 55;
			5165: Pixel = 114;
			5166: Pixel = 78;
			5167: Pixel = 45;
			5168: Pixel = 54;
			5169: Pixel = 46;
			5170: Pixel = 42;
			5171: Pixel = 117;
			5172: Pixel = 132;
			5173: Pixel = 65;
			5174: Pixel = 66;
			5175: Pixel = 49;
			5176: Pixel = 49;
			5177: Pixel = 50;
			5178: Pixel = 51;
			5179: Pixel = 124;
			5180: Pixel = 142;
			5181: Pixel = 155;
			5182: Pixel = 159;
			5183: Pixel = 155;
			5184: Pixel = 153;
			5185: Pixel = 153;
			5186: Pixel = 153;
			5187: Pixel = 153;
			5188: Pixel = 153;
			5189: Pixel = 154;
			5190: Pixel = 153;
			5191: Pixel = 153;
			5192: Pixel = 152;
			5193: Pixel = 149;
			5194: Pixel = 150;
			5195: Pixel = 145;
			5196: Pixel = 142;
			5197: Pixel = 137;
			5198: Pixel = 135;
			5199: Pixel = 131;
			5200: Pixel = 99;
			5201: Pixel = 97;
			5202: Pixel = 95;
			5203: Pixel = 88;
			5204: Pixel = 74;
			5205: Pixel = 100;
			5206: Pixel = 148;
			5207: Pixel = 171;
			5208: Pixel = 177;
			5209: Pixel = 179;
			5210: Pixel = 175;
			5211: Pixel = 150;
			5212: Pixel = 104;
			5213: Pixel = 76;
			5214: Pixel = 91;
			5215: Pixel = 100;
			5216: Pixel = 101;
			5217: Pixel = 100;
			5218: Pixel = 109;
			5219: Pixel = 84;
			5220: Pixel = 70;
			5221: Pixel = 136;
			5222: Pixel = 171;
			5223: Pixel = 177;
			5224: Pixel = 101;
			5225: Pixel = 60;
			5226: Pixel = 47;
			5227: Pixel = 82;
			5228: Pixel = 60;
			5229: Pixel = 64;
			5230: Pixel = 59;
			5231: Pixel = 107;
			5232: Pixel = 90;
			5233: Pixel = 41;
			5234: Pixel = 43;
			5235: Pixel = 58;
			5236: Pixel = 72;
			5237: Pixel = 40;
			5238: Pixel = 44;
			5239: Pixel = 42;
			5240: Pixel = 42;
			5241: Pixel = 91;
			5242: Pixel = 146;
			5243: Pixel = 169;
			5244: Pixel = 186;
			5245: Pixel = 206;
			5246: Pixel = 151;
			5247: Pixel = 102;
			5248: Pixel = 82;
			5249: Pixel = 56;
			5250: Pixel = 100;
			5251: Pixel = 72;
			5252: Pixel = 89;
			5253: Pixel = 206;
			5254: Pixel = 194;
			5255: Pixel = 103;
			5256: Pixel = 107;
			5257: Pixel = 118;
			5258: Pixel = 132;
			5259: Pixel = 152;
			5260: Pixel = 203;
			5261: Pixel = 195;
			5262: Pixel = 92;
			5263: Pixel = 75;
			5264: Pixel = 72;
			5265: Pixel = 151;
			5266: Pixel = 121;
			5267: Pixel = 40;
			5268: Pixel = 47;
			5269: Pixel = 45;
			5270: Pixel = 49;
			5271: Pixel = 113;
			5272: Pixel = 137;
			5273: Pixel = 75;
			5274: Pixel = 64;
			5275: Pixel = 49;
			5276: Pixel = 53;
			5277: Pixel = 44;
			5278: Pixel = 71;
			5279: Pixel = 140;
			5280: Pixel = 141;
			5281: Pixel = 157;
			5282: Pixel = 156;
			5283: Pixel = 155;
			5284: Pixel = 152;
			5285: Pixel = 152;
			5286: Pixel = 151;
			5287: Pixel = 153;
			5288: Pixel = 152;
			5289: Pixel = 152;
			5290: Pixel = 152;
			5291: Pixel = 150;
			5292: Pixel = 148;
			5293: Pixel = 146;
			5294: Pixel = 144;
			5295: Pixel = 140;
			5296: Pixel = 134;
			5297: Pixel = 127;
			5298: Pixel = 132;
			5299: Pixel = 146;
			5300: Pixel = 101;
			5301: Pixel = 99;
			5302: Pixel = 96;
			5303: Pixel = 89;
			5304: Pixel = 73;
			5305: Pixel = 98;
			5306: Pixel = 148;
			5307: Pixel = 169;
			5308: Pixel = 178;
			5309: Pixel = 180;
			5310: Pixel = 176;
			5311: Pixel = 152;
			5312: Pixel = 107;
			5313: Pixel = 82;
			5314: Pixel = 94;
			5315: Pixel = 104;
			5316: Pixel = 109;
			5317: Pixel = 108;
			5318: Pixel = 64;
			5319: Pixel = 74;
			5320: Pixel = 114;
			5321: Pixel = 162;
			5322: Pixel = 195;
			5323: Pixel = 122;
			5324: Pixel = 55;
			5325: Pixel = 50;
			5326: Pixel = 93;
			5327: Pixel = 60;
			5328: Pixel = 59;
			5329: Pixel = 79;
			5330: Pixel = 88;
			5331: Pixel = 110;
			5332: Pixel = 106;
			5333: Pixel = 56;
			5334: Pixel = 46;
			5335: Pixel = 44;
			5336: Pixel = 53;
			5337: Pixel = 49;
			5338: Pixel = 50;
			5339: Pixel = 31;
			5340: Pixel = 66;
			5341: Pixel = 132;
			5342: Pixel = 167;
			5343: Pixel = 180;
			5344: Pixel = 206;
			5345: Pixel = 148;
			5346: Pixel = 113;
			5347: Pixel = 133;
			5348: Pixel = 141;
			5349: Pixel = 102;
			5350: Pixel = 110;
			5351: Pixel = 117;
			5352: Pixel = 157;
			5353: Pixel = 193;
			5354: Pixel = 175;
			5355: Pixel = 139;
			5356: Pixel = 123;
			5357: Pixel = 121;
			5358: Pixel = 129;
			5359: Pixel = 153;
			5360: Pixel = 214;
			5361: Pixel = 179;
			5362: Pixel = 117;
			5363: Pixel = 127;
			5364: Pixel = 133;
			5365: Pixel = 162;
			5366: Pixel = 90;
			5367: Pixel = 53;
			5368: Pixel = 53;
			5369: Pixel = 49;
			5370: Pixel = 55;
			5371: Pixel = 105;
			5372: Pixel = 144;
			5373: Pixel = 79;
			5374: Pixel = 61;
			5375: Pixel = 46;
			5376: Pixel = 53;
			5377: Pixel = 46;
			5378: Pixel = 94;
			5379: Pixel = 141;
			5380: Pixel = 146;
			5381: Pixel = 158;
			5382: Pixel = 154;
			5383: Pixel = 152;
			5384: Pixel = 150;
			5385: Pixel = 153;
			5386: Pixel = 156;
			5387: Pixel = 152;
			5388: Pixel = 154;
			5389: Pixel = 152;
			5390: Pixel = 150;
			5391: Pixel = 147;
			5392: Pixel = 145;
			5393: Pixel = 142;
			5394: Pixel = 139;
			5395: Pixel = 132;
			5396: Pixel = 135;
			5397: Pixel = 152;
			5398: Pixel = 169;
			5399: Pixel = 183;
			5400: Pixel = 103;
			5401: Pixel = 102;
			5402: Pixel = 94;
			5403: Pixel = 86;
			5404: Pixel = 72;
			5405: Pixel = 97;
			5406: Pixel = 148;
			5407: Pixel = 170;
			5408: Pixel = 178;
			5409: Pixel = 182;
			5410: Pixel = 179;
			5411: Pixel = 155;
			5412: Pixel = 108;
			5413: Pixel = 81;
			5414: Pixel = 97;
			5415: Pixel = 107;
			5416: Pixel = 112;
			5417: Pixel = 115;
			5418: Pixel = 84;
			5419: Pixel = 145;
			5420: Pixel = 140;
			5421: Pixel = 125;
			5422: Pixel = 89;
			5423: Pixel = 30;
			5424: Pixel = 76;
			5425: Pixel = 111;
			5426: Pixel = 100;
			5427: Pixel = 50;
			5428: Pixel = 62;
			5429: Pixel = 84;
			5430: Pixel = 77;
			5431: Pixel = 112;
			5432: Pixel = 125;
			5433: Pixel = 80;
			5434: Pixel = 42;
			5435: Pixel = 46;
			5436: Pixel = 46;
			5437: Pixel = 49;
			5438: Pixel = 42;
			5439: Pixel = 37;
			5440: Pixel = 110;
			5441: Pixel = 154;
			5442: Pixel = 177;
			5443: Pixel = 204;
			5444: Pixel = 145;
			5445: Pixel = 103;
			5446: Pixel = 137;
			5447: Pixel = 141;
			5448: Pixel = 146;
			5449: Pixel = 145;
			5450: Pixel = 132;
			5451: Pixel = 121;
			5452: Pixel = 130;
			5453: Pixel = 130;
			5454: Pixel = 156;
			5455: Pixel = 157;
			5456: Pixel = 128;
			5457: Pixel = 128;
			5458: Pixel = 128;
			5459: Pixel = 147;
			5460: Pixel = 208;
			5461: Pixel = 202;
			5462: Pixel = 150;
			5463: Pixel = 135;
			5464: Pixel = 129;
			5465: Pixel = 96;
			5466: Pixel = 75;
			5467: Pixel = 82;
			5468: Pixel = 53;
			5469: Pixel = 49;
			5470: Pixel = 58;
			5471: Pixel = 95;
			5472: Pixel = 158;
			5473: Pixel = 80;
			5474: Pixel = 56;
			5475: Pixel = 47;
			5476: Pixel = 53;
			5477: Pixel = 56;
			5478: Pixel = 123;
			5479: Pixel = 137;
			5480: Pixel = 154;
			5481: Pixel = 156;
			5482: Pixel = 153;
			5483: Pixel = 152;
			5484: Pixel = 150;
			5485: Pixel = 151;
			5486: Pixel = 153;
			5487: Pixel = 150;
			5488: Pixel = 151;
			5489: Pixel = 151;
			5490: Pixel = 146;
			5491: Pixel = 142;
			5492: Pixel = 139;
			5493: Pixel = 134;
			5494: Pixel = 134;
			5495: Pixel = 151;
			5496: Pixel = 174;
			5497: Pixel = 187;
			5498: Pixel = 189;
			5499: Pixel = 188;
			5500: Pixel = 99;
			5501: Pixel = 95;
			5502: Pixel = 87;
			5503: Pixel = 83;
			5504: Pixel = 64;
			5505: Pixel = 89;
			5506: Pixel = 147;
			5507: Pixel = 169;
			5508: Pixel = 179;
			5509: Pixel = 182;
			5510: Pixel = 179;
			5511: Pixel = 156;
			5512: Pixel = 109;
			5513: Pixel = 79;
			5514: Pixel = 95;
			5515: Pixel = 106;
			5516: Pixel = 105;
			5517: Pixel = 112;
			5518: Pixel = 150;
			5519: Pixel = 132;
			5520: Pixel = 80;
			5521: Pixel = 76;
			5522: Pixel = 55;
			5523: Pixel = 53;
			5524: Pixel = 67;
			5525: Pixel = 103;
			5526: Pixel = 109;
			5527: Pixel = 62;
			5528: Pixel = 52;
			5529: Pixel = 76;
			5530: Pixel = 96;
			5531: Pixel = 96;
			5532: Pixel = 109;
			5533: Pixel = 76;
			5534: Pixel = 43;
			5535: Pixel = 46;
			5536: Pixel = 46;
			5537: Pixel = 51;
			5538: Pixel = 34;
			5539: Pixel = 81;
			5540: Pixel = 135;
			5541: Pixel = 169;
			5542: Pixel = 200;
			5543: Pixel = 155;
			5544: Pixel = 86;
			5545: Pixel = 123;
			5546: Pixel = 140;
			5547: Pixel = 152;
			5548: Pixel = 155;
			5549: Pixel = 156;
			5550: Pixel = 154;
			5551: Pixel = 150;
			5552: Pixel = 154;
			5553: Pixel = 163;
			5554: Pixel = 164;
			5555: Pixel = 156;
			5556: Pixel = 134;
			5557: Pixel = 136;
			5558: Pixel = 126;
			5559: Pixel = 142;
			5560: Pixel = 202;
			5561: Pixel = 209;
			5562: Pixel = 169;
			5563: Pixel = 149;
			5564: Pixel = 135;
			5565: Pixel = 120;
			5566: Pixel = 112;
			5567: Pixel = 96;
			5568: Pixel = 55;
			5569: Pixel = 49;
			5570: Pixel = 57;
			5571: Pixel = 89;
			5572: Pixel = 165;
			5573: Pixel = 78;
			5574: Pixel = 52;
			5575: Pixel = 48;
			5576: Pixel = 47;
			5577: Pixel = 63;
			5578: Pixel = 134;
			5579: Pixel = 138;
			5580: Pixel = 157;
			5581: Pixel = 154;
			5582: Pixel = 152;
			5583: Pixel = 150;
			5584: Pixel = 151;
			5585: Pixel = 151;
			5586: Pixel = 149;
			5587: Pixel = 150;
			5588: Pixel = 149;
			5589: Pixel = 147;
			5590: Pixel = 144;
			5591: Pixel = 142;
			5592: Pixel = 134;
			5593: Pixel = 133;
			5594: Pixel = 166;
			5595: Pixel = 190;
			5596: Pixel = 193;
			5597: Pixel = 191;
			5598: Pixel = 189;
			5599: Pixel = 189;
			5600: Pixel = 94;
			5601: Pixel = 89;
			5602: Pixel = 83;
			5603: Pixel = 78;
			5604: Pixel = 60;
			5605: Pixel = 87;
			5606: Pixel = 145;
			5607: Pixel = 168;
			5608: Pixel = 178;
			5609: Pixel = 181;
			5610: Pixel = 178;
			5611: Pixel = 156;
			5612: Pixel = 109;
			5613: Pixel = 80;
			5614: Pixel = 93;
			5615: Pixel = 103;
			5616: Pixel = 115;
			5617: Pixel = 124;
			5618: Pixel = 135;
			5619: Pixel = 126;
			5620: Pixel = 112;
			5621: Pixel = 80;
			5622: Pixel = 52;
			5623: Pixel = 80;
			5624: Pixel = 106;
			5625: Pixel = 99;
			5626: Pixel = 81;
			5627: Pixel = 38;
			5628: Pixel = 53;
			5629: Pixel = 87;
			5630: Pixel = 97;
			5631: Pixel = 113;
			5632: Pixel = 112;
			5633: Pixel = 84;
			5634: Pixel = 56;
			5635: Pixel = 47;
			5636: Pixel = 46;
			5637: Pixel = 46;
			5638: Pixel = 54;
			5639: Pixel = 118;
			5640: Pixel = 148;
			5641: Pixel = 200;
			5642: Pixel = 171;
			5643: Pixel = 69;
			5644: Pixel = 109;
			5645: Pixel = 127;
			5646: Pixel = 138;
			5647: Pixel = 151;
			5648: Pixel = 162;
			5649: Pixel = 168;
			5650: Pixel = 173;
			5651: Pixel = 170;
			5652: Pixel = 173;
			5653: Pixel = 172;
			5654: Pixel = 171;
			5655: Pixel = 154;
			5656: Pixel = 141;
			5657: Pixel = 137;
			5658: Pixel = 126;
			5659: Pixel = 136;
			5660: Pixel = 195;
			5661: Pixel = 213;
			5662: Pixel = 177;
			5663: Pixel = 160;
			5664: Pixel = 142;
			5665: Pixel = 132;
			5666: Pixel = 125;
			5667: Pixel = 105;
			5668: Pixel = 58;
			5669: Pixel = 54;
			5670: Pixel = 56;
			5671: Pixel = 78;
			5672: Pixel = 172;
			5673: Pixel = 77;
			5674: Pixel = 46;
			5675: Pixel = 50;
			5676: Pixel = 42;
			5677: Pixel = 87;
			5678: Pixel = 138;
			5679: Pixel = 145;
			5680: Pixel = 158;
			5681: Pixel = 153;
			5682: Pixel = 152;
			5683: Pixel = 151;
			5684: Pixel = 150;
			5685: Pixel = 151;
			5686: Pixel = 148;
			5687: Pixel = 147;
			5688: Pixel = 146;
			5689: Pixel = 143;
			5690: Pixel = 141;
			5691: Pixel = 136;
			5692: Pixel = 134;
			5693: Pixel = 169;
			5694: Pixel = 197;
			5695: Pixel = 197;
			5696: Pixel = 192;
			5697: Pixel = 189;
			5698: Pixel = 188;
			5699: Pixel = 190;
			5700: Pixel = 88;
			5701: Pixel = 84;
			5702: Pixel = 80;
			5703: Pixel = 75;
			5704: Pixel = 58;
			5705: Pixel = 87;
			5706: Pixel = 145;
			5707: Pixel = 169;
			5708: Pixel = 177;
			5709: Pixel = 181;
			5710: Pixel = 178;
			5711: Pixel = 156;
			5712: Pixel = 108;
			5713: Pixel = 78;
			5714: Pixel = 92;
			5715: Pixel = 112;
			5716: Pixel = 129;
			5717: Pixel = 136;
			5718: Pixel = 119;
			5719: Pixel = 85;
			5720: Pixel = 73;
			5721: Pixel = 54;
			5722: Pixel = 75;
			5723: Pixel = 89;
			5724: Pixel = 113;
			5725: Pixel = 107;
			5726: Pixel = 57;
			5727: Pixel = 44;
			5728: Pixel = 43;
			5729: Pixel = 59;
			5730: Pixel = 88;
			5731: Pixel = 82;
			5732: Pixel = 52;
			5733: Pixel = 126;
			5734: Pixel = 83;
			5735: Pixel = 42;
			5736: Pixel = 48;
			5737: Pixel = 36;
			5738: Pixel = 91;
			5739: Pixel = 133;
			5740: Pixel = 180;
			5741: Pixel = 196;
			5742: Pixel = 65;
			5743: Pixel = 74;
			5744: Pixel = 120;
			5745: Pixel = 124;
			5746: Pixel = 136;
			5747: Pixel = 148;
			5748: Pixel = 159;
			5749: Pixel = 171;
			5750: Pixel = 176;
			5751: Pixel = 177;
			5752: Pixel = 175;
			5753: Pixel = 175;
			5754: Pixel = 170;
			5755: Pixel = 155;
			5756: Pixel = 147;
			5757: Pixel = 139;
			5758: Pixel = 129;
			5759: Pixel = 132;
			5760: Pixel = 188;
			5761: Pixel = 218;
			5762: Pixel = 174;
			5763: Pixel = 160;
			5764: Pixel = 144;
			5765: Pixel = 132;
			5766: Pixel = 129;
			5767: Pixel = 107;
			5768: Pixel = 56;
			5769: Pixel = 58;
			5770: Pixel = 60;
			5771: Pixel = 68;
			5772: Pixel = 168;
			5773: Pixel = 86;
			5774: Pixel = 38;
			5775: Pixel = 52;
			5776: Pixel = 43;
			5777: Pixel = 111;
			5778: Pixel = 141;
			5779: Pixel = 152;
			5780: Pixel = 158;
			5781: Pixel = 153;
			5782: Pixel = 152;
			5783: Pixel = 151;
			5784: Pixel = 150;
			5785: Pixel = 150;
			5786: Pixel = 148;
			5787: Pixel = 145;
			5788: Pixel = 145;
			5789: Pixel = 142;
			5790: Pixel = 136;
			5791: Pixel = 130;
			5792: Pixel = 163;
			5793: Pixel = 194;
			5794: Pixel = 195;
			5795: Pixel = 195;
			5796: Pixel = 193;
			5797: Pixel = 190;
			5798: Pixel = 193;
			5799: Pixel = 198;
			5800: Pixel = 79;
			5801: Pixel = 76;
			5802: Pixel = 74;
			5803: Pixel = 72;
			5804: Pixel = 57;
			5805: Pixel = 84;
			5806: Pixel = 144;
			5807: Pixel = 168;
			5808: Pixel = 176;
			5809: Pixel = 178;
			5810: Pixel = 175;
			5811: Pixel = 155;
			5812: Pixel = 109;
			5813: Pixel = 78;
			5814: Pixel = 92;
			5815: Pixel = 105;
			5816: Pixel = 109;
			5817: Pixel = 106;
			5818: Pixel = 98;
			5819: Pixel = 92;
			5820: Pixel = 83;
			5821: Pixel = 83;
			5822: Pixel = 79;
			5823: Pixel = 76;
			5824: Pixel = 116;
			5825: Pixel = 69;
			5826: Pixel = 50;
			5827: Pixel = 49;
			5828: Pixel = 51;
			5829: Pixel = 49;
			5830: Pixel = 55;
			5831: Pixel = 51;
			5832: Pixel = 46;
			5833: Pixel = 120;
			5834: Pixel = 117;
			5835: Pixel = 38;
			5836: Pixel = 36;
			5837: Pixel = 48;
			5838: Pixel = 119;
			5839: Pixel = 155;
			5840: Pixel = 210;
			5841: Pixel = 105;
			5842: Pixel = 35;
			5843: Pixel = 91;
			5844: Pixel = 121;
			5845: Pixel = 126;
			5846: Pixel = 134;
			5847: Pixel = 144;
			5848: Pixel = 152;
			5849: Pixel = 164;
			5850: Pixel = 174;
			5851: Pixel = 179;
			5852: Pixel = 176;
			5853: Pixel = 172;
			5854: Pixel = 164;
			5855: Pixel = 150;
			5856: Pixel = 144;
			5857: Pixel = 139;
			5858: Pixel = 127;
			5859: Pixel = 133;
			5860: Pixel = 180;
			5861: Pixel = 220;
			5862: Pixel = 176;
			5863: Pixel = 158;
			5864: Pixel = 149;
			5865: Pixel = 135;
			5866: Pixel = 130;
			5867: Pixel = 100;
			5868: Pixel = 51;
			5869: Pixel = 54;
			5870: Pixel = 61;
			5871: Pixel = 59;
			5872: Pixel = 165;
			5873: Pixel = 102;
			5874: Pixel = 37;
			5875: Pixel = 56;
			5876: Pixel = 54;
			5877: Pixel = 127;
			5878: Pixel = 145;
			5879: Pixel = 162;
			5880: Pixel = 155;
			5881: Pixel = 153;
			5882: Pixel = 152;
			5883: Pixel = 149;
			5884: Pixel = 148;
			5885: Pixel = 147;
			5886: Pixel = 146;
			5887: Pixel = 145;
			5888: Pixel = 144;
			5889: Pixel = 140;
			5890: Pixel = 129;
			5891: Pixel = 146;
			5892: Pixel = 190;
			5893: Pixel = 195;
			5894: Pixel = 192;
			5895: Pixel = 193;
			5896: Pixel = 194;
			5897: Pixel = 197;
			5898: Pixel = 203;
			5899: Pixel = 204;
			5900: Pixel = 76;
			5901: Pixel = 75;
			5902: Pixel = 74;
			5903: Pixel = 68;
			5904: Pixel = 52;
			5905: Pixel = 83;
			5906: Pixel = 144;
			5907: Pixel = 166;
			5908: Pixel = 173;
			5909: Pixel = 174;
			5910: Pixel = 174;
			5911: Pixel = 154;
			5912: Pixel = 108;
			5913: Pixel = 75;
			5914: Pixel = 107;
			5915: Pixel = 101;
			5916: Pixel = 126;
			5917: Pixel = 124;
			5918: Pixel = 88;
			5919: Pixel = 105;
			5920: Pixel = 103;
			5921: Pixel = 78;
			5922: Pixel = 67;
			5923: Pixel = 73;
			5924: Pixel = 120;
			5925: Pixel = 80;
			5926: Pixel = 55;
			5927: Pixel = 56;
			5928: Pixel = 44;
			5929: Pixel = 42;
			5930: Pixel = 66;
			5931: Pixel = 55;
			5932: Pixel = 65;
			5933: Pixel = 117;
			5934: Pixel = 123;
			5935: Pixel = 98;
			5936: Pixel = 22;
			5937: Pixel = 84;
			5938: Pixel = 126;
			5939: Pixel = 200;
			5940: Pixel = 166;
			5941: Pixel = 35;
			5942: Pixel = 57;
			5943: Pixel = 84;
			5944: Pixel = 117;
			5945: Pixel = 127;
			5946: Pixel = 134;
			5947: Pixel = 143;
			5948: Pixel = 152;
			5949: Pixel = 157;
			5950: Pixel = 168;
			5951: Pixel = 174;
			5952: Pixel = 173;
			5953: Pixel = 169;
			5954: Pixel = 161;
			5955: Pixel = 145;
			5956: Pixel = 135;
			5957: Pixel = 133;
			5958: Pixel = 124;
			5959: Pixel = 131;
			5960: Pixel = 168;
			5961: Pixel = 220;
			5962: Pixel = 178;
			5963: Pixel = 154;
			5964: Pixel = 148;
			5965: Pixel = 135;
			5966: Pixel = 129;
			5967: Pixel = 88;
			5968: Pixel = 45;
			5969: Pixel = 59;
			5970: Pixel = 63;
			5971: Pixel = 51;
			5972: Pixel = 158;
			5973: Pixel = 119;
			5974: Pixel = 43;
			5975: Pixel = 49;
			5976: Pixel = 75;
			5977: Pixel = 138;
			5978: Pixel = 149;
			5979: Pixel = 163;
			5980: Pixel = 155;
			5981: Pixel = 154;
			5982: Pixel = 152;
			5983: Pixel = 149;
			5984: Pixel = 147;
			5985: Pixel = 145;
			5986: Pixel = 144;
			5987: Pixel = 143;
			5988: Pixel = 141;
			5989: Pixel = 135;
			5990: Pixel = 132;
			5991: Pixel = 176;
			5992: Pixel = 197;
			5993: Pixel = 192;
			5994: Pixel = 192;
			5995: Pixel = 195;
			5996: Pixel = 201;
			5997: Pixel = 207;
			5998: Pixel = 205;
			5999: Pixel = 202;
			6000: Pixel = 78;
			6001: Pixel = 76;
			6002: Pixel = 74;
			6003: Pixel = 66;
			6004: Pixel = 49;
			6005: Pixel = 81;
			6006: Pixel = 143;
			6007: Pixel = 166;
			6008: Pixel = 172;
			6009: Pixel = 174;
			6010: Pixel = 173;
			6011: Pixel = 154;
			6012: Pixel = 107;
			6013: Pixel = 70;
			6014: Pixel = 107;
			6015: Pixel = 126;
			6016: Pixel = 135;
			6017: Pixel = 101;
			6018: Pixel = 71;
			6019: Pixel = 114;
			6020: Pixel = 86;
			6021: Pixel = 64;
			6022: Pixel = 97;
			6023: Pixel = 99;
			6024: Pixel = 125;
			6025: Pixel = 97;
			6026: Pixel = 53;
			6027: Pixel = 53;
			6028: Pixel = 37;
			6029: Pixel = 46;
			6030: Pixel = 89;
			6031: Pixel = 73;
			6032: Pixel = 96;
			6033: Pixel = 163;
			6034: Pixel = 88;
			6035: Pixel = 70;
			6036: Pixel = 31;
			6037: Pixel = 114;
			6038: Pixel = 157;
			6039: Pixel = 199;
			6040: Pixel = 57;
			6041: Pixel = 36;
			6042: Pixel = 67;
			6043: Pixel = 80;
			6044: Pixel = 114;
			6045: Pixel = 127;
			6046: Pixel = 131;
			6047: Pixel = 139;
			6048: Pixel = 149;
			6049: Pixel = 156;
			6050: Pixel = 159;
			6051: Pixel = 164;
			6052: Pixel = 167;
			6053: Pixel = 165;
			6054: Pixel = 159;
			6055: Pixel = 141;
			6056: Pixel = 131;
			6057: Pixel = 128;
			6058: Pixel = 120;
			6059: Pixel = 126;
			6060: Pixel = 159;
			6061: Pixel = 217;
			6062: Pixel = 188;
			6063: Pixel = 150;
			6064: Pixel = 147;
			6065: Pixel = 135;
			6066: Pixel = 125;
			6067: Pixel = 71;
			6068: Pixel = 42;
			6069: Pixel = 66;
			6070: Pixel = 66;
			6071: Pixel = 43;
			6072: Pixel = 148;
			6073: Pixel = 131;
			6074: Pixel = 43;
			6075: Pixel = 42;
			6076: Pixel = 98;
			6077: Pixel = 143;
			6078: Pixel = 152;
			6079: Pixel = 159;
			6080: Pixel = 153;
			6081: Pixel = 153;
			6082: Pixel = 153;
			6083: Pixel = 150;
			6084: Pixel = 147;
			6085: Pixel = 147;
			6086: Pixel = 145;
			6087: Pixel = 141;
			6088: Pixel = 139;
			6089: Pixel = 130;
			6090: Pixel = 154;
			6091: Pixel = 194;
			6092: Pixel = 194;
			6093: Pixel = 192;
			6094: Pixel = 194;
			6095: Pixel = 203;
			6096: Pixel = 207;
			6097: Pixel = 208;
			6098: Pixel = 205;
			6099: Pixel = 203;
			6100: Pixel = 81;
			6101: Pixel = 77;
			6102: Pixel = 74;
			6103: Pixel = 63;
			6104: Pixel = 43;
			6105: Pixel = 75;
			6106: Pixel = 142;
			6107: Pixel = 167;
			6108: Pixel = 174;
			6109: Pixel = 176;
			6110: Pixel = 176;
			6111: Pixel = 156;
			6112: Pixel = 107;
			6113: Pixel = 70;
			6114: Pixel = 98;
			6115: Pixel = 117;
			6116: Pixel = 120;
			6117: Pixel = 96;
			6118: Pixel = 78;
			6119: Pixel = 95;
			6120: Pixel = 84;
			6121: Pixel = 80;
			6122: Pixel = 92;
			6123: Pixel = 83;
			6124: Pixel = 122;
			6125: Pixel = 92;
			6126: Pixel = 47;
			6127: Pixel = 50;
			6128: Pixel = 46;
			6129: Pixel = 51;
			6130: Pixel = 82;
			6131: Pixel = 110;
			6132: Pixel = 111;
			6133: Pixel = 86;
			6134: Pixel = 54;
			6135: Pixel = 32;
			6136: Pixel = 87;
			6137: Pixel = 116;
			6138: Pixel = 180;
			6139: Pixel = 111;
			6140: Pixel = 23;
			6141: Pixel = 49;
			6142: Pixel = 78;
			6143: Pixel = 79;
			6144: Pixel = 112;
			6145: Pixel = 125;
			6146: Pixel = 131;
			6147: Pixel = 137;
			6148: Pixel = 145;
			6149: Pixel = 151;
			6150: Pixel = 152;
			6151: Pixel = 157;
			6152: Pixel = 161;
			6153: Pixel = 161;
			6154: Pixel = 152;
			6155: Pixel = 132;
			6156: Pixel = 121;
			6157: Pixel = 137;
			6158: Pixel = 131;
			6159: Pixel = 126;
			6160: Pixel = 152;
			6161: Pixel = 215;
			6162: Pixel = 197;
			6163: Pixel = 144;
			6164: Pixel = 146;
			6165: Pixel = 133;
			6166: Pixel = 116;
			6167: Pixel = 52;
			6168: Pixel = 45;
			6169: Pixel = 67;
			6170: Pixel = 65;
			6171: Pixel = 37;
			6172: Pixel = 134;
			6173: Pixel = 149;
			6174: Pixel = 52;
			6175: Pixel = 43;
			6176: Pixel = 124;
			6177: Pixel = 144;
			6178: Pixel = 156;
			6179: Pixel = 156;
			6180: Pixel = 152;
			6181: Pixel = 150;
			6182: Pixel = 150;
			6183: Pixel = 150;
			6184: Pixel = 149;
			6185: Pixel = 147;
			6186: Pixel = 146;
			6187: Pixel = 143;
			6188: Pixel = 135;
			6189: Pixel = 134;
			6190: Pixel = 181;
			6191: Pixel = 198;
			6192: Pixel = 193;
			6193: Pixel = 194;
			6194: Pixel = 202;
			6195: Pixel = 208;
			6196: Pixel = 205;
			6197: Pixel = 205;
			6198: Pixel = 207;
			6199: Pixel = 207;
			6200: Pixel = 84;
			6201: Pixel = 80;
			6202: Pixel = 74;
			6203: Pixel = 66;
			6204: Pixel = 45;
			6205: Pixel = 78;
			6206: Pixel = 142;
			6207: Pixel = 167;
			6208: Pixel = 173;
			6209: Pixel = 176;
			6210: Pixel = 177;
			6211: Pixel = 156;
			6212: Pixel = 110;
			6213: Pixel = 90;
			6214: Pixel = 112;
			6215: Pixel = 103;
			6216: Pixel = 117;
			6217: Pixel = 80;
			6218: Pixel = 81;
			6219: Pixel = 112;
			6220: Pixel = 67;
			6221: Pixel = 84;
			6222: Pixel = 79;
			6223: Pixel = 75;
			6224: Pixel = 118;
			6225: Pixel = 101;
			6226: Pixel = 71;
			6227: Pixel = 53;
			6228: Pixel = 53;
			6229: Pixel = 41;
			6230: Pixel = 78;
			6231: Pixel = 69;
			6232: Pixel = 99;
			6233: Pixel = 46;
			6234: Pixel = 24;
			6235: Pixel = 75;
			6236: Pixel = 175;
			6237: Pixel = 160;
			6238: Pixel = 156;
			6239: Pixel = 54;
			6240: Pixel = 36;
			6241: Pixel = 49;
			6242: Pixel = 85;
			6243: Pixel = 81;
			6244: Pixel = 114;
			6245: Pixel = 125;
			6246: Pixel = 129;
			6247: Pixel = 137;
			6248: Pixel = 143;
			6249: Pixel = 148;
			6250: Pixel = 151;
			6251: Pixel = 154;
			6252: Pixel = 158;
			6253: Pixel = 158;
			6254: Pixel = 152;
			6255: Pixel = 127;
			6256: Pixel = 125;
			6257: Pixel = 128;
			6258: Pixel = 125;
			6259: Pixel = 123;
			6260: Pixel = 142;
			6261: Pixel = 203;
			6262: Pixel = 183;
			6263: Pixel = 142;
			6264: Pixel = 142;
			6265: Pixel = 132;
			6266: Pixel = 89;
			6267: Pixel = 39;
			6268: Pixel = 49;
			6269: Pixel = 66;
			6270: Pixel = 64;
			6271: Pixel = 34;
			6272: Pixel = 119;
			6273: Pixel = 160;
			6274: Pixel = 60;
			6275: Pixel = 51;
			6276: Pixel = 142;
			6277: Pixel = 148;
			6278: Pixel = 158;
			6279: Pixel = 154;
			6280: Pixel = 151;
			6281: Pixel = 149;
			6282: Pixel = 149;
			6283: Pixel = 149;
			6284: Pixel = 148;
			6285: Pixel = 147;
			6286: Pixel = 145;
			6287: Pixel = 142;
			6288: Pixel = 130;
			6289: Pixel = 150;
			6290: Pixel = 194;
			6291: Pixel = 195;
			6292: Pixel = 193;
			6293: Pixel = 199;
			6294: Pixel = 206;
			6295: Pixel = 206;
			6296: Pixel = 205;
			6297: Pixel = 206;
			6298: Pixel = 208;
			6299: Pixel = 207;
			6300: Pixel = 80;
			6301: Pixel = 78;
			6302: Pixel = 76;
			6303: Pixel = 68;
			6304: Pixel = 59;
			6305: Pixel = 96;
			6306: Pixel = 148;
			6307: Pixel = 166;
			6308: Pixel = 172;
			6309: Pixel = 175;
			6310: Pixel = 177;
			6311: Pixel = 157;
			6312: Pixel = 114;
			6313: Pixel = 78;
			6314: Pixel = 87;
			6315: Pixel = 103;
			6316: Pixel = 111;
			6317: Pixel = 82;
			6318: Pixel = 88;
			6319: Pixel = 102;
			6320: Pixel = 54;
			6321: Pixel = 105;
			6322: Pixel = 76;
			6323: Pixel = 77;
			6324: Pixel = 115;
			6325: Pixel = 123;
			6326: Pixel = 82;
			6327: Pixel = 42;
			6328: Pixel = 76;
			6329: Pixel = 50;
			6330: Pixel = 31;
			6331: Pixel = 93;
			6332: Pixel = 73;
			6333: Pixel = 41;
			6334: Pixel = 38;
			6335: Pixel = 115;
			6336: Pixel = 181;
			6337: Pixel = 185;
			6338: Pixel = 65;
			6339: Pixel = 35;
			6340: Pixel = 44;
			6341: Pixel = 49;
			6342: Pixel = 92;
			6343: Pixel = 91;
			6344: Pixel = 113;
			6345: Pixel = 123;
			6346: Pixel = 129;
			6347: Pixel = 135;
			6348: Pixel = 142;
			6349: Pixel = 148;
			6350: Pixel = 150;
			6351: Pixel = 152;
			6352: Pixel = 156;
			6353: Pixel = 158;
			6354: Pixel = 153;
			6355: Pixel = 138;
			6356: Pixel = 127;
			6357: Pixel = 104;
			6358: Pixel = 98;
			6359: Pixel = 105;
			6360: Pixel = 121;
			6361: Pixel = 177;
			6362: Pixel = 166;
			6363: Pixel = 145;
			6364: Pixel = 139;
			6365: Pixel = 125;
			6366: Pixel = 58;
			6367: Pixel = 43;
			6368: Pixel = 53;
			6369: Pixel = 69;
			6370: Pixel = 63;
			6371: Pixel = 36;
			6372: Pixel = 100;
			6373: Pixel = 163;
			6374: Pixel = 69;
			6375: Pixel = 79;
			6376: Pixel = 150;
			6377: Pixel = 150;
			6378: Pixel = 158;
			6379: Pixel = 152;
			6380: Pixel = 150;
			6381: Pixel = 149;
			6382: Pixel = 150;
			6383: Pixel = 148;
			6384: Pixel = 146;
			6385: Pixel = 144;
			6386: Pixel = 144;
			6387: Pixel = 141;
			6388: Pixel = 131;
			6389: Pixel = 166;
			6390: Pixel = 197;
			6391: Pixel = 195;
			6392: Pixel = 198;
			6393: Pixel = 206;
			6394: Pixel = 206;
			6395: Pixel = 206;
			6396: Pixel = 209;
			6397: Pixel = 209;
			6398: Pixel = 209;
			6399: Pixel = 206;
			6400: Pixel = 79;
			6401: Pixel = 77;
			6402: Pixel = 76;
			6403: Pixel = 69;
			6404: Pixel = 73;
			6405: Pixel = 111;
			6406: Pixel = 153;
			6407: Pixel = 166;
			6408: Pixel = 169;
			6409: Pixel = 174;
			6410: Pixel = 178;
			6411: Pixel = 159;
			6412: Pixel = 112;
			6413: Pixel = 75;
			6414: Pixel = 91;
			6415: Pixel = 102;
			6416: Pixel = 120;
			6417: Pixel = 69;
			6418: Pixel = 74;
			6419: Pixel = 61;
			6420: Pixel = 87;
			6421: Pixel = 79;
			6422: Pixel = 75;
			6423: Pixel = 94;
			6424: Pixel = 104;
			6425: Pixel = 124;
			6426: Pixel = 116;
			6427: Pixel = 34;
			6428: Pixel = 93;
			6429: Pixel = 110;
			6430: Pixel = 34;
			6431: Pixel = 76;
			6432: Pixel = 65;
			6433: Pixel = 102;
			6434: Pixel = 137;
			6435: Pixel = 106;
			6436: Pixel = 162;
			6437: Pixel = 103;
			6438: Pixel = 30;
			6439: Pixel = 63;
			6440: Pixel = 48;
			6441: Pixel = 50;
			6442: Pixel = 100;
			6443: Pixel = 94;
			6444: Pixel = 117;
			6445: Pixel = 123;
			6446: Pixel = 127;
			6447: Pixel = 132;
			6448: Pixel = 140;
			6449: Pixel = 145;
			6450: Pixel = 146;
			6451: Pixel = 151;
			6452: Pixel = 154;
			6453: Pixel = 158;
			6454: Pixel = 156;
			6455: Pixel = 151;
			6456: Pixel = 139;
			6457: Pixel = 134;
			6458: Pixel = 143;
			6459: Pixel = 139;
			6460: Pixel = 174;
			6461: Pixel = 186;
			6462: Pixel = 159;
			6463: Pixel = 144;
			6464: Pixel = 138;
			6465: Pixel = 98;
			6466: Pixel = 43;
			6467: Pixel = 48;
			6468: Pixel = 57;
			6469: Pixel = 78;
			6470: Pixel = 68;
			6471: Pixel = 41;
			6472: Pixel = 83;
			6473: Pixel = 160;
			6474: Pixel = 79;
			6475: Pixel = 105;
			6476: Pixel = 152;
			6477: Pixel = 153;
			6478: Pixel = 156;
			6479: Pixel = 152;
			6480: Pixel = 151;
			6481: Pixel = 149;
			6482: Pixel = 148;
			6483: Pixel = 148;
			6484: Pixel = 146;
			6485: Pixel = 145;
			6486: Pixel = 143;
			6487: Pixel = 137;
			6488: Pixel = 134;
			6489: Pixel = 179;
			6490: Pixel = 197;
			6491: Pixel = 196;
			6492: Pixel = 204;
			6493: Pixel = 207;
			6494: Pixel = 206;
			6495: Pixel = 207;
			6496: Pixel = 210;
			6497: Pixel = 209;
			6498: Pixel = 207;
			6499: Pixel = 208;
			6500: Pixel = 75;
			6501: Pixel = 75;
			6502: Pixel = 77;
			6503: Pixel = 65;
			6504: Pixel = 72;
			6505: Pixel = 120;
			6506: Pixel = 154;
			6507: Pixel = 165;
			6508: Pixel = 169;
			6509: Pixel = 176;
			6510: Pixel = 178;
			6511: Pixel = 159;
			6512: Pixel = 114;
			6513: Pixel = 76;
			6514: Pixel = 87;
			6515: Pixel = 104;
			6516: Pixel = 136;
			6517: Pixel = 70;
			6518: Pixel = 70;
			6519: Pixel = 101;
			6520: Pixel = 77;
			6521: Pixel = 48;
			6522: Pixel = 72;
			6523: Pixel = 88;
			6524: Pixel = 102;
			6525: Pixel = 101;
			6526: Pixel = 133;
			6527: Pixel = 78;
			6528: Pixel = 84;
			6529: Pixel = 85;
			6530: Pixel = 44;
			6531: Pixel = 72;
			6532: Pixel = 139;
			6533: Pixel = 174;
			6534: Pixel = 127;
			6535: Pixel = 114;
			6536: Pixel = 141;
			6537: Pixel = 40;
			6538: Pixel = 52;
			6539: Pixel = 57;
			6540: Pixel = 56;
			6541: Pixel = 50;
			6542: Pixel = 99;
			6543: Pixel = 99;
			6544: Pixel = 118;
			6545: Pixel = 125;
			6546: Pixel = 127;
			6547: Pixel = 134;
			6548: Pixel = 140;
			6549: Pixel = 141;
			6550: Pixel = 143;
			6551: Pixel = 150;
			6552: Pixel = 153;
			6553: Pixel = 155;
			6554: Pixel = 155;
			6555: Pixel = 151;
			6556: Pixel = 149;
			6557: Pixel = 143;
			6558: Pixel = 176;
			6559: Pixel = 182;
			6560: Pixel = 194;
			6561: Pixel = 189;
			6562: Pixel = 154;
			6563: Pixel = 142;
			6564: Pixel = 133;
			6565: Pixel = 64;
			6566: Pixel = 45;
			6567: Pixel = 48;
			6568: Pixel = 65;
			6569: Pixel = 78;
			6570: Pixel = 68;
			6571: Pixel = 48;
			6572: Pixel = 66;
			6573: Pixel = 154;
			6574: Pixel = 96;
			6575: Pixel = 127;
			6576: Pixel = 149;
			6577: Pixel = 155;
			6578: Pixel = 154;
			6579: Pixel = 151;
			6580: Pixel = 150;
			6581: Pixel = 148;
			6582: Pixel = 147;
			6583: Pixel = 145;
			6584: Pixel = 146;
			6585: Pixel = 145;
			6586: Pixel = 142;
			6587: Pixel = 135;
			6588: Pixel = 140;
			6589: Pixel = 186;
			6590: Pixel = 196;
			6591: Pixel = 200;
			6592: Pixel = 208;
			6593: Pixel = 207;
			6594: Pixel = 205;
			6595: Pixel = 207;
			6596: Pixel = 208;
			6597: Pixel = 210;
			6598: Pixel = 210;
			6599: Pixel = 211;
			6600: Pixel = 72;
			6601: Pixel = 70;
			6602: Pixel = 70;
			6603: Pixel = 63;
			6604: Pixel = 73;
			6605: Pixel = 117;
			6606: Pixel = 153;
			6607: Pixel = 166;
			6608: Pixel = 170;
			6609: Pixel = 175;
			6610: Pixel = 178;
			6611: Pixel = 161;
			6612: Pixel = 114;
			6613: Pixel = 73;
			6614: Pixel = 86;
			6615: Pixel = 123;
			6616: Pixel = 118;
			6617: Pixel = 72;
			6618: Pixel = 101;
			6619: Pixel = 79;
			6620: Pixel = 55;
			6621: Pixel = 67;
			6622: Pixel = 69;
			6623: Pixel = 68;
			6624: Pixel = 85;
			6625: Pixel = 80;
			6626: Pixel = 123;
			6627: Pixel = 119;
			6628: Pixel = 90;
			6629: Pixel = 44;
			6630: Pixel = 73;
			6631: Pixel = 107;
			6632: Pixel = 170;
			6633: Pixel = 167;
			6634: Pixel = 90;
			6635: Pixel = 130;
			6636: Pixel = 51;
			6637: Pixel = 49;
			6638: Pixel = 49;
			6639: Pixel = 56;
			6640: Pixel = 62;
			6641: Pixel = 43;
			6642: Pixel = 94;
			6643: Pixel = 99;
			6644: Pixel = 113;
			6645: Pixel = 126;
			6646: Pixel = 128;
			6647: Pixel = 133;
			6648: Pixel = 140;
			6649: Pixel = 140;
			6650: Pixel = 139;
			6651: Pixel = 142;
			6652: Pixel = 148;
			6653: Pixel = 148;
			6654: Pixel = 150;
			6655: Pixel = 147;
			6656: Pixel = 150;
			6657: Pixel = 156;
			6658: Pixel = 196;
			6659: Pixel = 196;
			6660: Pixel = 199;
			6661: Pixel = 193;
			6662: Pixel = 149;
			6663: Pixel = 144;
			6664: Pixel = 107;
			6665: Pixel = 42;
			6666: Pixel = 50;
			6667: Pixel = 50;
			6668: Pixel = 68;
			6669: Pixel = 76;
			6670: Pixel = 66;
			6671: Pixel = 48;
			6672: Pixel = 56;
			6673: Pixel = 145;
			6674: Pixel = 110;
			6675: Pixel = 137;
			6676: Pixel = 149;
			6677: Pixel = 155;
			6678: Pixel = 153;
			6679: Pixel = 151;
			6680: Pixel = 148;
			6681: Pixel = 148;
			6682: Pixel = 147;
			6683: Pixel = 145;
			6684: Pixel = 145;
			6685: Pixel = 144;
			6686: Pixel = 142;
			6687: Pixel = 131;
			6688: Pixel = 145;
			6689: Pixel = 191;
			6690: Pixel = 198;
			6691: Pixel = 206;
			6692: Pixel = 208;
			6693: Pixel = 207;
			6694: Pixel = 208;
			6695: Pixel = 206;
			6696: Pixel = 209;
			6697: Pixel = 211;
			6698: Pixel = 210;
			6699: Pixel = 211;
			6700: Pixel = 65;
			6701: Pixel = 64;
			6702: Pixel = 69;
			6703: Pixel = 64;
			6704: Pixel = 71;
			6705: Pixel = 113;
			6706: Pixel = 154;
			6707: Pixel = 167;
			6708: Pixel = 171;
			6709: Pixel = 176;
			6710: Pixel = 179;
			6711: Pixel = 162;
			6712: Pixel = 114;
			6713: Pixel = 67;
			6714: Pixel = 110;
			6715: Pixel = 108;
			6716: Pixel = 112;
			6717: Pixel = 64;
			6718: Pixel = 91;
			6719: Pixel = 66;
			6720: Pixel = 61;
			6721: Pixel = 64;
			6722: Pixel = 82;
			6723: Pixel = 85;
			6724: Pixel = 76;
			6725: Pixel = 77;
			6726: Pixel = 79;
			6727: Pixel = 133;
			6728: Pixel = 79;
			6729: Pixel = 72;
			6730: Pixel = 151;
			6731: Pixel = 171;
			6732: Pixel = 180;
			6733: Pixel = 98;
			6734: Pixel = 128;
			6735: Pixel = 73;
			6736: Pixel = 44;
			6737: Pixel = 70;
			6738: Pixel = 44;
			6739: Pixel = 59;
			6740: Pixel = 69;
			6741: Pixel = 43;
			6742: Pixel = 87;
			6743: Pixel = 91;
			6744: Pixel = 106;
			6745: Pixel = 125;
			6746: Pixel = 129;
			6747: Pixel = 132;
			6748: Pixel = 137;
			6749: Pixel = 140;
			6750: Pixel = 137;
			6751: Pixel = 138;
			6752: Pixel = 132;
			6753: Pixel = 138;
			6754: Pixel = 143;
			6755: Pixel = 142;
			6756: Pixel = 145;
			6757: Pixel = 147;
			6758: Pixel = 155;
			6759: Pixel = 173;
			6760: Pixel = 164;
			6761: Pixel = 156;
			6762: Pixel = 130;
			6763: Pixel = 141;
			6764: Pixel = 68;
			6765: Pixel = 43;
			6766: Pixel = 53;
			6767: Pixel = 52;
			6768: Pixel = 69;
			6769: Pixel = 77;
			6770: Pixel = 71;
			6771: Pixel = 51;
			6772: Pixel = 47;
			6773: Pixel = 140;
			6774: Pixel = 122;
			6775: Pixel = 141;
			6776: Pixel = 148;
			6777: Pixel = 156;
			6778: Pixel = 152;
			6779: Pixel = 150;
			6780: Pixel = 147;
			6781: Pixel = 148;
			6782: Pixel = 148;
			6783: Pixel = 146;
			6784: Pixel = 145;
			6785: Pixel = 144;
			6786: Pixel = 141;
			6787: Pixel = 129;
			6788: Pixel = 148;
			6789: Pixel = 193;
			6790: Pixel = 203;
			6791: Pixel = 209;
			6792: Pixel = 208;
			6793: Pixel = 208;
			6794: Pixel = 209;
			6795: Pixel = 208;
			6796: Pixel = 211;
			6797: Pixel = 212;
			6798: Pixel = 211;
			6799: Pixel = 212;
			6800: Pixel = 56;
			6801: Pixel = 59;
			6802: Pixel = 65;
			6803: Pixel = 62;
			6804: Pixel = 74;
			6805: Pixel = 117;
			6806: Pixel = 156;
			6807: Pixel = 170;
			6808: Pixel = 175;
			6809: Pixel = 178;
			6810: Pixel = 179;
			6811: Pixel = 160;
			6812: Pixel = 106;
			6813: Pixel = 97;
			6814: Pixel = 108;
			6815: Pixel = 104;
			6816: Pixel = 128;
			6817: Pixel = 58;
			6818: Pixel = 60;
			6819: Pixel = 63;
			6820: Pixel = 68;
			6821: Pixel = 53;
			6822: Pixel = 95;
			6823: Pixel = 115;
			6824: Pixel = 93;
			6825: Pixel = 80;
			6826: Pixel = 101;
			6827: Pixel = 87;
			6828: Pixel = 90;
			6829: Pixel = 129;
			6830: Pixel = 167;
			6831: Pixel = 221;
			6832: Pixel = 113;
			6833: Pixel = 115;
			6834: Pixel = 118;
			6835: Pixel = 35;
			6836: Pixel = 51;
			6837: Pixel = 58;
			6838: Pixel = 45;
			6839: Pixel = 57;
			6840: Pixel = 69;
			6841: Pixel = 46;
			6842: Pixel = 80;
			6843: Pixel = 84;
			6844: Pixel = 98;
			6845: Pixel = 123;
			6846: Pixel = 128;
			6847: Pixel = 127;
			6848: Pixel = 134;
			6849: Pixel = 139;
			6850: Pixel = 145;
			6851: Pixel = 134;
			6852: Pixel = 100;
			6853: Pixel = 102;
			6854: Pixel = 110;
			6855: Pixel = 116;
			6856: Pixel = 110;
			6857: Pixel = 101;
			6858: Pixel = 109;
			6859: Pixel = 126;
			6860: Pixel = 107;
			6861: Pixel = 110;
			6862: Pixel = 134;
			6863: Pixel = 117;
			6864: Pixel = 41;
			6865: Pixel = 51;
			6866: Pixel = 47;
			6867: Pixel = 58;
			6868: Pixel = 67;
			6869: Pixel = 77;
			6870: Pixel = 66;
			6871: Pixel = 59;
			6872: Pixel = 44;
			6873: Pixel = 127;
			6874: Pixel = 140;
			6875: Pixel = 146;
			6876: Pixel = 150;
			6877: Pixel = 156;
			6878: Pixel = 152;
			6879: Pixel = 151;
			6880: Pixel = 149;
			6881: Pixel = 147;
			6882: Pixel = 147;
			6883: Pixel = 146;
			6884: Pixel = 144;
			6885: Pixel = 144;
			6886: Pixel = 141;
			6887: Pixel = 127;
			6888: Pixel = 153;
			6889: Pixel = 198;
			6890: Pixel = 209;
			6891: Pixel = 210;
			6892: Pixel = 209;
			6893: Pixel = 208;
			6894: Pixel = 209;
			6895: Pixel = 210;
			6896: Pixel = 211;
			6897: Pixel = 213;
			6898: Pixel = 213;
			6899: Pixel = 213;
			6900: Pixel = 56;
			6901: Pixel = 59;
			6902: Pixel = 63;
			6903: Pixel = 62;
			6904: Pixel = 83;
			6905: Pixel = 119;
			6906: Pixel = 154;
			6907: Pixel = 170;
			6908: Pixel = 176;
			6909: Pixel = 180;
			6910: Pixel = 179;
			6911: Pixel = 157;
			6912: Pixel = 127;
			6913: Pixel = 113;
			6914: Pixel = 79;
			6915: Pixel = 129;
			6916: Pixel = 109;
			6917: Pixel = 70;
			6918: Pixel = 65;
			6919: Pixel = 44;
			6920: Pixel = 69;
			6921: Pixel = 63;
			6922: Pixel = 112;
			6923: Pixel = 103;
			6924: Pixel = 88;
			6925: Pixel = 105;
			6926: Pixel = 84;
			6927: Pixel = 80;
			6928: Pixel = 113;
			6929: Pixel = 135;
			6930: Pixel = 161;
			6931: Pixel = 162;
			6932: Pixel = 109;
			6933: Pixel = 149;
			6934: Pixel = 52;
			6935: Pixel = 50;
			6936: Pixel = 45;
			6937: Pixel = 53;
			6938: Pixel = 49;
			6939: Pixel = 56;
			6940: Pixel = 65;
			6941: Pixel = 53;
			6942: Pixel = 71;
			6943: Pixel = 79;
			6944: Pixel = 91;
			6945: Pixel = 116;
			6946: Pixel = 121;
			6947: Pixel = 124;
			6948: Pixel = 129;
			6949: Pixel = 135;
			6950: Pixel = 145;
			6951: Pixel = 145;
			6952: Pixel = 133;
			6953: Pixel = 121;
			6954: Pixel = 119;
			6955: Pixel = 125;
			6956: Pixel = 139;
			6957: Pixel = 158;
			6958: Pixel = 167;
			6959: Pixel = 181;
			6960: Pixel = 147;
			6961: Pixel = 142;
			6962: Pixel = 144;
			6963: Pixel = 62;
			6964: Pixel = 43;
			6965: Pixel = 50;
			6966: Pixel = 47;
			6967: Pixel = 55;
			6968: Pixel = 67;
			6969: Pixel = 80;
			6970: Pixel = 65;
			6971: Pixel = 69;
			6972: Pixel = 44;
			6973: Pixel = 122;
			6974: Pixel = 153;
			6975: Pixel = 147;
			6976: Pixel = 152;
			6977: Pixel = 155;
			6978: Pixel = 152;
			6979: Pixel = 152;
			6980: Pixel = 151;
			6981: Pixel = 148;
			6982: Pixel = 147;
			6983: Pixel = 146;
			6984: Pixel = 145;
			6985: Pixel = 145;
			6986: Pixel = 140;
			6987: Pixel = 125;
			6988: Pixel = 159;
			6989: Pixel = 207;
			6990: Pixel = 212;
			6991: Pixel = 210;
			6992: Pixel = 210;
			6993: Pixel = 210;
			6994: Pixel = 211;
			6995: Pixel = 212;
			6996: Pixel = 213;
			6997: Pixel = 212;
			6998: Pixel = 211;
			6999: Pixel = 210;
			7000: Pixel = 54;
			7001: Pixel = 55;
			7002: Pixel = 58;
			7003: Pixel = 58;
			7004: Pixel = 82;
			7005: Pixel = 114;
			7006: Pixel = 153;
			7007: Pixel = 168;
			7008: Pixel = 177;
			7009: Pixel = 180;
			7010: Pixel = 178;
			7011: Pixel = 166;
			7012: Pixel = 125;
			7013: Pixel = 64;
			7014: Pixel = 104;
			7015: Pixel = 127;
			7016: Pixel = 84;
			7017: Pixel = 86;
			7018: Pixel = 82;
			7019: Pixel = 42;
			7020: Pixel = 79;
			7021: Pixel = 73;
			7022: Pixel = 126;
			7023: Pixel = 106;
			7024: Pixel = 78;
			7025: Pixel = 93;
			7026: Pixel = 101;
			7027: Pixel = 101;
			7028: Pixel = 145;
			7029: Pixel = 137;
			7030: Pixel = 157;
			7031: Pixel = 135;
			7032: Pixel = 167;
			7033: Pixel = 71;
			7034: Pixel = 46;
			7035: Pixel = 57;
			7036: Pixel = 49;
			7037: Pixel = 51;
			7038: Pixel = 51;
			7039: Pixel = 56;
			7040: Pixel = 66;
			7041: Pixel = 56;
			7042: Pixel = 69;
			7043: Pixel = 74;
			7044: Pixel = 78;
			7045: Pixel = 106;
			7046: Pixel = 113;
			7047: Pixel = 119;
			7048: Pixel = 125;
			7049: Pixel = 131;
			7050: Pixel = 138;
			7051: Pixel = 144;
			7052: Pixel = 141;
			7053: Pixel = 131;
			7054: Pixel = 127;
			7055: Pixel = 125;
			7056: Pixel = 130;
			7057: Pixel = 146;
			7058: Pixel = 146;
			7059: Pixel = 141;
			7060: Pixel = 142;
			7061: Pixel = 151;
			7062: Pixel = 101;
			7063: Pixel = 39;
			7064: Pixel = 50;
			7065: Pixel = 49;
			7066: Pixel = 51;
			7067: Pixel = 52;
			7068: Pixel = 68;
			7069: Pixel = 81;
			7070: Pixel = 70;
			7071: Pixel = 70;
			7072: Pixel = 47;
			7073: Pixel = 122;
			7074: Pixel = 159;
			7075: Pixel = 149;
			7076: Pixel = 153;
			7077: Pixel = 155;
			7078: Pixel = 153;
			7079: Pixel = 153;
			7080: Pixel = 152;
			7081: Pixel = 150;
			7082: Pixel = 149;
			7083: Pixel = 146;
			7084: Pixel = 144;
			7085: Pixel = 143;
			7086: Pixel = 139;
			7087: Pixel = 123;
			7088: Pixel = 164;
			7089: Pixel = 214;
			7090: Pixel = 214;
			7091: Pixel = 211;
			7092: Pixel = 211;
			7093: Pixel = 214;
			7094: Pixel = 214;
			7095: Pixel = 213;
			7096: Pixel = 210;
			7097: Pixel = 206;
			7098: Pixel = 205;
			7099: Pixel = 204;
			7100: Pixel = 51;
			7101: Pixel = 52;
			7102: Pixel = 51;
			7103: Pixel = 59;
			7104: Pixel = 89;
			7105: Pixel = 108;
			7106: Pixel = 147;
			7107: Pixel = 166;
			7108: Pixel = 178;
			7109: Pixel = 179;
			7110: Pixel = 179;
			7111: Pixel = 160;
			7112: Pixel = 107;
			7113: Pixel = 66;
			7114: Pixel = 122;
			7115: Pixel = 107;
			7116: Pixel = 65;
			7117: Pixel = 90;
			7118: Pixel = 67;
			7119: Pixel = 52;
			7120: Pixel = 70;
			7121: Pixel = 66;
			7122: Pixel = 144;
			7123: Pixel = 104;
			7124: Pixel = 122;
			7125: Pixel = 80;
			7126: Pixel = 113;
			7127: Pixel = 121;
			7128: Pixel = 108;
			7129: Pixel = 128;
			7130: Pixel = 168;
			7131: Pixel = 183;
			7132: Pixel = 91;
			7133: Pixel = 41;
			7134: Pixel = 55;
			7135: Pixel = 57;
			7136: Pixel = 52;
			7137: Pixel = 52;
			7138: Pixel = 55;
			7139: Pixel = 60;
			7140: Pixel = 62;
			7141: Pixel = 58;
			7142: Pixel = 62;
			7143: Pixel = 72;
			7144: Pixel = 68;
			7145: Pixel = 92;
			7146: Pixel = 104;
			7147: Pixel = 112;
			7148: Pixel = 122;
			7149: Pixel = 129;
			7150: Pixel = 134;
			7151: Pixel = 139;
			7152: Pixel = 139;
			7153: Pixel = 135;
			7154: Pixel = 130;
			7155: Pixel = 129;
			7156: Pixel = 125;
			7157: Pixel = 124;
			7158: Pixel = 128;
			7159: Pixel = 140;
			7160: Pixel = 149;
			7161: Pixel = 125;
			7162: Pixel = 59;
			7163: Pixel = 43;
			7164: Pixel = 47;
			7165: Pixel = 56;
			7166: Pixel = 57;
			7167: Pixel = 50;
			7168: Pixel = 73;
			7169: Pixel = 83;
			7170: Pixel = 70;
			7171: Pixel = 71;
			7172: Pixel = 50;
			7173: Pixel = 118;
			7174: Pixel = 162;
			7175: Pixel = 148;
			7176: Pixel = 154;
			7177: Pixel = 154;
			7178: Pixel = 153;
			7179: Pixel = 154;
			7180: Pixel = 154;
			7181: Pixel = 153;
			7182: Pixel = 149;
			7183: Pixel = 147;
			7184: Pixel = 143;
			7185: Pixel = 141;
			7186: Pixel = 136;
			7187: Pixel = 118;
			7188: Pixel = 165;
			7189: Pixel = 219;
			7190: Pixel = 215;
			7191: Pixel = 213;
			7192: Pixel = 214;
			7193: Pixel = 217;
			7194: Pixel = 213;
			7195: Pixel = 208;
			7196: Pixel = 205;
			7197: Pixel = 206;
			7198: Pixel = 208;
			7199: Pixel = 209;
			7200: Pixel = 50;
			7201: Pixel = 51;
			7202: Pixel = 45;
			7203: Pixel = 69;
			7204: Pixel = 103;
			7205: Pixel = 114;
			7206: Pixel = 142;
			7207: Pixel = 164;
			7208: Pixel = 176;
			7209: Pixel = 177;
			7210: Pixel = 178;
			7211: Pixel = 160;
			7212: Pixel = 114;
			7213: Pixel = 68;
			7214: Pixel = 110;
			7215: Pixel = 99;
			7216: Pixel = 73;
			7217: Pixel = 83;
			7218: Pixel = 48;
			7219: Pixel = 58;
			7220: Pixel = 64;
			7221: Pixel = 63;
			7222: Pixel = 134;
			7223: Pixel = 113;
			7224: Pixel = 131;
			7225: Pixel = 113;
			7226: Pixel = 89;
			7227: Pixel = 111;
			7228: Pixel = 98;
			7229: Pixel = 111;
			7230: Pixel = 196;
			7231: Pixel = 120;
			7232: Pixel = 37;
			7233: Pixel = 54;
			7234: Pixel = 50;
			7235: Pixel = 57;
			7236: Pixel = 50;
			7237: Pixel = 53;
			7238: Pixel = 51;
			7239: Pixel = 52;
			7240: Pixel = 58;
			7241: Pixel = 59;
			7242: Pixel = 52;
			7243: Pixel = 64;
			7244: Pixel = 61;
			7245: Pixel = 73;
			7246: Pixel = 93;
			7247: Pixel = 106;
			7248: Pixel = 118;
			7249: Pixel = 128;
			7250: Pixel = 133;
			7251: Pixel = 137;
			7252: Pixel = 138;
			7253: Pixel = 140;
			7254: Pixel = 143;
			7255: Pixel = 146;
			7256: Pixel = 159;
			7257: Pixel = 163;
			7258: Pixel = 157;
			7259: Pixel = 154;
			7260: Pixel = 149;
			7261: Pixel = 81;
			7262: Pixel = 48;
			7263: Pixel = 45;
			7264: Pixel = 51;
			7265: Pixel = 60;
			7266: Pixel = 56;
			7267: Pixel = 47;
			7268: Pixel = 79;
			7269: Pixel = 84;
			7270: Pixel = 74;
			7271: Pixel = 76;
			7272: Pixel = 51;
			7273: Pixel = 115;
			7274: Pixel = 166;
			7275: Pixel = 147;
			7276: Pixel = 156;
			7277: Pixel = 155;
			7278: Pixel = 154;
			7279: Pixel = 153;
			7280: Pixel = 152;
			7281: Pixel = 152;
			7282: Pixel = 149;
			7283: Pixel = 147;
			7284: Pixel = 143;
			7285: Pixel = 141;
			7286: Pixel = 133;
			7287: Pixel = 115;
			7288: Pixel = 167;
			7289: Pixel = 221;
			7290: Pixel = 216;
			7291: Pixel = 214;
			7292: Pixel = 214;
			7293: Pixel = 213;
			7294: Pixel = 211;
			7295: Pixel = 211;
			7296: Pixel = 211;
			7297: Pixel = 209;
			7298: Pixel = 208;
			7299: Pixel = 207;
			7300: Pixel = 47;
			7301: Pixel = 49;
			7302: Pixel = 46;
			7303: Pixel = 74;
			7304: Pixel = 101;
			7305: Pixel = 114;
			7306: Pixel = 143;
			7307: Pixel = 165;
			7308: Pixel = 176;
			7309: Pixel = 176;
			7310: Pixel = 177;
			7311: Pixel = 160;
			7312: Pixel = 112;
			7313: Pixel = 69;
			7314: Pixel = 96;
			7315: Pixel = 92;
			7316: Pixel = 69;
			7317: Pixel = 86;
			7318: Pixel = 48;
			7319: Pixel = 62;
			7320: Pixel = 58;
			7321: Pixel = 67;
			7322: Pixel = 109;
			7323: Pixel = 77;
			7324: Pixel = 111;
			7325: Pixel = 131;
			7326: Pixel = 100;
			7327: Pixel = 111;
			7328: Pixel = 127;
			7329: Pixel = 91;
			7330: Pixel = 130;
			7331: Pixel = 63;
			7332: Pixel = 50;
			7333: Pixel = 51;
			7334: Pixel = 53;
			7335: Pixel = 60;
			7336: Pixel = 49;
			7337: Pixel = 53;
			7338: Pixel = 51;
			7339: Pixel = 47;
			7340: Pixel = 54;
			7341: Pixel = 57;
			7342: Pixel = 54;
			7343: Pixel = 59;
			7344: Pixel = 60;
			7345: Pixel = 63;
			7346: Pixel = 59;
			7347: Pixel = 87;
			7348: Pixel = 105;
			7349: Pixel = 126;
			7350: Pixel = 134;
			7351: Pixel = 137;
			7352: Pixel = 143;
			7353: Pixel = 147;
			7354: Pixel = 161;
			7355: Pixel = 163;
			7356: Pixel = 167;
			7357: Pixel = 169;
			7358: Pixel = 168;
			7359: Pixel = 157;
			7360: Pixel = 135;
			7361: Pixel = 54;
			7362: Pixel = 53;
			7363: Pixel = 47;
			7364: Pixel = 56;
			7365: Pixel = 59;
			7366: Pixel = 55;
			7367: Pixel = 50;
			7368: Pixel = 86;
			7369: Pixel = 87;
			7370: Pixel = 76;
			7371: Pixel = 75;
			7372: Pixel = 55;
			7373: Pixel = 114;
			7374: Pixel = 168;
			7375: Pixel = 147;
			7376: Pixel = 158;
			7377: Pixel = 155;
			7378: Pixel = 151;
			7379: Pixel = 150;
			7380: Pixel = 149;
			7381: Pixel = 151;
			7382: Pixel = 149;
			7383: Pixel = 146;
			7384: Pixel = 140;
			7385: Pixel = 138;
			7386: Pixel = 132;
			7387: Pixel = 116;
			7388: Pixel = 180;
			7389: Pixel = 223;
			7390: Pixel = 215;
			7391: Pixel = 211;
			7392: Pixel = 212;
			7393: Pixel = 213;
			7394: Pixel = 213;
			7395: Pixel = 209;
			7396: Pixel = 206;
			7397: Pixel = 206;
			7398: Pixel = 211;
			7399: Pixel = 210;
			7400: Pixel = 48;
			7401: Pixel = 48;
			7402: Pixel = 45;
			7403: Pixel = 63;
			7404: Pixel = 94;
			7405: Pixel = 120;
			7406: Pixel = 144;
			7407: Pixel = 166;
			7408: Pixel = 174;
			7409: Pixel = 176;
			7410: Pixel = 178;
			7411: Pixel = 162;
			7412: Pixel = 113;
			7413: Pixel = 58;
			7414: Pixel = 96;
			7415: Pixel = 65;
			7416: Pixel = 57;
			7417: Pixel = 86;
			7418: Pixel = 55;
			7419: Pixel = 65;
			7420: Pixel = 54;
			7421: Pixel = 56;
			7422: Pixel = 127;
			7423: Pixel = 66;
			7424: Pixel = 78;
			7425: Pixel = 116;
			7426: Pixel = 131;
			7427: Pixel = 125;
			7428: Pixel = 138;
			7429: Pixel = 108;
			7430: Pixel = 77;
			7431: Pixel = 53;
			7432: Pixel = 54;
			7433: Pixel = 51;
			7434: Pixel = 54;
			7435: Pixel = 63;
			7436: Pixel = 51;
			7437: Pixel = 56;
			7438: Pixel = 53;
			7439: Pixel = 51;
			7440: Pixel = 49;
			7441: Pixel = 56;
			7442: Pixel = 57;
			7443: Pixel = 59;
			7444: Pixel = 59;
			7445: Pixel = 69;
			7446: Pixel = 52;
			7447: Pixel = 50;
			7448: Pixel = 74;
			7449: Pixel = 99;
			7450: Pixel = 112;
			7451: Pixel = 125;
			7452: Pixel = 136;
			7453: Pixel = 144;
			7454: Pixel = 152;
			7455: Pixel = 163;
			7456: Pixel = 168;
			7457: Pixel = 163;
			7458: Pixel = 162;
			7459: Pixel = 153;
			7460: Pixel = 110;
			7461: Pixel = 48;
			7462: Pixel = 59;
			7463: Pixel = 55;
			7464: Pixel = 57;
			7465: Pixel = 61;
			7466: Pixel = 52;
			7467: Pixel = 53;
			7468: Pixel = 90;
			7469: Pixel = 86;
			7470: Pixel = 79;
			7471: Pixel = 81;
			7472: Pixel = 60;
			7473: Pixel = 114;
			7474: Pixel = 168;
			7475: Pixel = 143;
			7476: Pixel = 150;
			7477: Pixel = 151;
			7478: Pixel = 149;
			7479: Pixel = 151;
			7480: Pixel = 150;
			7481: Pixel = 149;
			7482: Pixel = 147;
			7483: Pixel = 142;
			7484: Pixel = 139;
			7485: Pixel = 137;
			7486: Pixel = 128;
			7487: Pixel = 119;
			7488: Pixel = 193;
			7489: Pixel = 224;
			7490: Pixel = 212;
			7491: Pixel = 210;
			7492: Pixel = 213;
			7493: Pixel = 214;
			7494: Pixel = 211;
			7495: Pixel = 206;
			7496: Pixel = 208;
			7497: Pixel = 200;
			7498: Pixel = 168;
			7499: Pixel = 125;
			7500: Pixel = 46;
			7501: Pixel = 46;
			7502: Pixel = 42;
			7503: Pixel = 53;
			7504: Pixel = 88;
			7505: Pixel = 111;
			7506: Pixel = 146;
			7507: Pixel = 167;
			7508: Pixel = 172;
			7509: Pixel = 174;
			7510: Pixel = 176;
			7511: Pixel = 160;
			7512: Pixel = 96;
			7513: Pixel = 103;
			7514: Pixel = 130;
			7515: Pixel = 80;
			7516: Pixel = 57;
			7517: Pixel = 73;
			7518: Pixel = 60;
			7519: Pixel = 62;
			7520: Pixel = 47;
			7521: Pixel = 44;
			7522: Pixel = 129;
			7523: Pixel = 114;
			7524: Pixel = 68;
			7525: Pixel = 101;
			7526: Pixel = 105;
			7527: Pixel = 114;
			7528: Pixel = 146;
			7529: Pixel = 131;
			7530: Pixel = 137;
			7531: Pixel = 71;
			7532: Pixel = 40;
			7533: Pixel = 51;
			7534: Pixel = 60;
			7535: Pixel = 70;
			7536: Pixel = 48;
			7537: Pixel = 58;
			7538: Pixel = 49;
			7539: Pixel = 52;
			7540: Pixel = 48;
			7541: Pixel = 51;
			7542: Pixel = 59;
			7543: Pixel = 62;
			7544: Pixel = 59;
			7545: Pixel = 63;
			7546: Pixel = 74;
			7547: Pixel = 62;
			7548: Pixel = 76;
			7549: Pixel = 86;
			7550: Pixel = 102;
			7551: Pixel = 114;
			7552: Pixel = 124;
			7553: Pixel = 135;
			7554: Pixel = 148;
			7555: Pixel = 155;
			7556: Pixel = 164;
			7557: Pixel = 161;
			7558: Pixel = 153;
			7559: Pixel = 148;
			7560: Pixel = 109;
			7561: Pixel = 45;
			7562: Pixel = 49;
			7563: Pixel = 55;
			7564: Pixel = 59;
			7565: Pixel = 61;
			7566: Pixel = 51;
			7567: Pixel = 55;
			7568: Pixel = 90;
			7569: Pixel = 90;
			7570: Pixel = 82;
			7571: Pixel = 83;
			7572: Pixel = 62;
			7573: Pixel = 123;
			7574: Pixel = 161;
			7575: Pixel = 119;
			7576: Pixel = 120;
			7577: Pixel = 132;
			7578: Pixel = 138;
			7579: Pixel = 142;
			7580: Pixel = 146;
			7581: Pixel = 149;
			7582: Pixel = 147;
			7583: Pixel = 143;
			7584: Pixel = 138;
			7585: Pixel = 134;
			7586: Pixel = 121;
			7587: Pixel = 130;
			7588: Pixel = 207;
			7589: Pixel = 218;
			7590: Pixel = 211;
			7591: Pixel = 210;
			7592: Pixel = 210;
			7593: Pixel = 210;
			7594: Pixel = 204;
			7595: Pixel = 195;
			7596: Pixel = 157;
			7597: Pixel = 93;
			7598: Pixel = 45;
			7599: Pixel = 38;
			7600: Pixel = 53;
			7601: Pixel = 52;
			7602: Pixel = 41;
			7603: Pixel = 48;
			7604: Pixel = 74;
			7605: Pixel = 97;
			7606: Pixel = 144;
			7607: Pixel = 165;
			7608: Pixel = 173;
			7609: Pixel = 172;
			7610: Pixel = 174;
			7611: Pixel = 148;
			7612: Pixel = 142;
			7613: Pixel = 139;
			7614: Pixel = 82;
			7615: Pixel = 79;
			7616: Pixel = 47;
			7617: Pixel = 78;
			7618: Pixel = 62;
			7619: Pixel = 63;
			7620: Pixel = 57;
			7621: Pixel = 47;
			7622: Pixel = 115;
			7623: Pixel = 134;
			7624: Pixel = 82;
			7625: Pixel = 62;
			7626: Pixel = 119;
			7627: Pixel = 113;
			7628: Pixel = 118;
			7629: Pixel = 120;
			7630: Pixel = 87;
			7631: Pixel = 152;
			7632: Pixel = 76;
			7633: Pixel = 39;
			7634: Pixel = 65;
			7635: Pixel = 70;
			7636: Pixel = 49;
			7637: Pixel = 59;
			7638: Pixel = 48;
			7639: Pixel = 52;
			7640: Pixel = 49;
			7641: Pixel = 50;
			7642: Pixel = 55;
			7643: Pixel = 59;
			7644: Pixel = 55;
			7645: Pixel = 52;
			7646: Pixel = 77;
			7647: Pixel = 100;
			7648: Pixel = 125;
			7649: Pixel = 130;
			7650: Pixel = 135;
			7651: Pixel = 137;
			7652: Pixel = 137;
			7653: Pixel = 142;
			7654: Pixel = 151;
			7655: Pixel = 153;
			7656: Pixel = 151;
			7657: Pixel = 155;
			7658: Pixel = 164;
			7659: Pixel = 182;
			7660: Pixel = 189;
			7661: Pixel = 160;
			7662: Pixel = 103;
			7663: Pixel = 56;
			7664: Pixel = 44;
			7665: Pixel = 54;
			7666: Pixel = 51;
			7667: Pixel = 57;
			7668: Pixel = 90;
			7669: Pixel = 89;
			7670: Pixel = 82;
			7671: Pixel = 84;
			7672: Pixel = 66;
			7673: Pixel = 131;
			7674: Pixel = 147;
			7675: Pixel = 112;
			7676: Pixel = 112;
			7677: Pixel = 113;
			7678: Pixel = 115;
			7679: Pixel = 117;
			7680: Pixel = 121;
			7681: Pixel = 129;
			7682: Pixel = 136;
			7683: Pixel = 137;
			7684: Pixel = 137;
			7685: Pixel = 133;
			7686: Pixel = 116;
			7687: Pixel = 146;
			7688: Pixel = 216;
			7689: Pixel = 210;
			7690: Pixel = 207;
			7691: Pixel = 209;
			7692: Pixel = 207;
			7693: Pixel = 202;
			7694: Pixel = 196;
			7695: Pixel = 148;
			7696: Pixel = 57;
			7697: Pixel = 33;
			7698: Pixel = 55;
			7699: Pixel = 73;
			7700: Pixel = 91;
			7701: Pixel = 70;
			7702: Pixel = 52;
			7703: Pixel = 53;
			7704: Pixel = 60;
			7705: Pixel = 76;
			7706: Pixel = 131;
			7707: Pixel = 164;
			7708: Pixel = 171;
			7709: Pixel = 170;
			7710: Pixel = 173;
			7711: Pixel = 173;
			7712: Pixel = 138;
			7713: Pixel = 61;
			7714: Pixel = 104;
			7715: Pixel = 57;
			7716: Pixel = 39;
			7717: Pixel = 72;
			7718: Pixel = 58;
			7719: Pixel = 57;
			7720: Pixel = 86;
			7721: Pixel = 59;
			7722: Pixel = 70;
			7723: Pixel = 122;
			7724: Pixel = 103;
			7725: Pixel = 100;
			7726: Pixel = 139;
			7727: Pixel = 88;
			7728: Pixel = 97;
			7729: Pixel = 111;
			7730: Pixel = 99;
			7731: Pixel = 136;
			7732: Pixel = 123;
			7733: Pixel = 61;
			7734: Pixel = 58;
			7735: Pixel = 65;
			7736: Pixel = 52;
			7737: Pixel = 63;
			7738: Pixel = 48;
			7739: Pixel = 50;
			7740: Pixel = 52;
			7741: Pixel = 49;
			7742: Pixel = 52;
			7743: Pixel = 60;
			7744: Pixel = 57;
			7745: Pixel = 52;
			7746: Pixel = 75;
			7747: Pixel = 110;
			7748: Pixel = 125;
			7749: Pixel = 124;
			7750: Pixel = 124;
			7751: Pixel = 132;
			7752: Pixel = 136;
			7753: Pixel = 139;
			7754: Pixel = 144;
			7755: Pixel = 141;
			7756: Pixel = 141;
			7757: Pixel = 146;
			7758: Pixel = 166;
			7759: Pixel = 185;
			7760: Pixel = 198;
			7761: Pixel = 208;
			7762: Pixel = 208;
			7763: Pixel = 177;
			7764: Pixel = 110;
			7765: Pixel = 48;
			7766: Pixel = 35;
			7767: Pixel = 56;
			7768: Pixel = 91;
			7769: Pixel = 84;
			7770: Pixel = 79;
			7771: Pixel = 80;
			7772: Pixel = 67;
			7773: Pixel = 135;
			7774: Pixel = 142;
			7775: Pixel = 128;
			7776: Pixel = 132;
			7777: Pixel = 123;
			7778: Pixel = 117;
			7779: Pixel = 109;
			7780: Pixel = 104;
			7781: Pixel = 102;
			7782: Pixel = 106;
			7783: Pixel = 111;
			7784: Pixel = 112;
			7785: Pixel = 116;
			7786: Pixel = 103;
			7787: Pixel = 146;
			7788: Pixel = 212;
			7789: Pixel = 204;
			7790: Pixel = 206;
			7791: Pixel = 208;
			7792: Pixel = 208;
			7793: Pixel = 199;
			7794: Pixel = 147;
			7795: Pixel = 65;
			7796: Pixel = 45;
			7797: Pixel = 64;
			7798: Pixel = 82;
			7799: Pixel = 86;
			7800: Pixel = 135;
			7801: Pixel = 117;
			7802: Pixel = 83;
			7803: Pixel = 71;
			7804: Pixel = 56;
			7805: Pixel = 60;
			7806: Pixel = 122;
			7807: Pixel = 163;
			7808: Pixel = 170;
			7809: Pixel = 170;
			7810: Pixel = 177;
			7811: Pixel = 167;
			7812: Pixel = 100;
			7813: Pixel = 120;
			7814: Pixel = 106;
			7815: Pixel = 33;
			7816: Pixel = 39;
			7817: Pixel = 67;
			7818: Pixel = 82;
			7819: Pixel = 34;
			7820: Pixel = 99;
			7821: Pixel = 89;
			7822: Pixel = 42;
			7823: Pixel = 83;
			7824: Pixel = 108;
			7825: Pixel = 110;
			7826: Pixel = 94;
			7827: Pixel = 92;
			7828: Pixel = 109;
			7829: Pixel = 116;
			7830: Pixel = 124;
			7831: Pixel = 130;
			7832: Pixel = 79;
			7833: Pixel = 102;
			7834: Pixel = 57;
			7835: Pixel = 59;
			7836: Pixel = 50;
			7837: Pixel = 63;
			7838: Pixel = 48;
			7839: Pixel = 48;
			7840: Pixel = 57;
			7841: Pixel = 51;
			7842: Pixel = 51;
			7843: Pixel = 59;
			7844: Pixel = 66;
			7845: Pixel = 52;
			7846: Pixel = 69;
			7847: Pixel = 107;
			7848: Pixel = 118;
			7849: Pixel = 123;
			7850: Pixel = 127;
			7851: Pixel = 130;
			7852: Pixel = 137;
			7853: Pixel = 139;
			7854: Pixel = 139;
			7855: Pixel = 139;
			7856: Pixel = 144;
			7857: Pixel = 154;
			7858: Pixel = 172;
			7859: Pixel = 187;
			7860: Pixel = 191;
			7861: Pixel = 193;
			7862: Pixel = 198;
			7863: Pixel = 208;
			7864: Pixel = 216;
			7865: Pixel = 173;
			7866: Pixel = 65;
			7867: Pixel = 38;
			7868: Pixel = 85;
			7869: Pixel = 80;
			7870: Pixel = 74;
			7871: Pixel = 74;
			7872: Pixel = 65;
			7873: Pixel = 137;
			7874: Pixel = 145;
			7875: Pixel = 141;
			7876: Pixel = 141;
			7877: Pixel = 136;
			7878: Pixel = 132;
			7879: Pixel = 127;
			7880: Pixel = 117;
			7881: Pixel = 108;
			7882: Pixel = 100;
			7883: Pixel = 93;
			7884: Pixel = 93;
			7885: Pixel = 117;
			7886: Pixel = 85;
			7887: Pixel = 124;
			7888: Pixel = 210;
			7889: Pixel = 205;
			7890: Pixel = 209;
			7891: Pixel = 207;
			7892: Pixel = 200;
			7893: Pixel = 150;
			7894: Pixel = 56;
			7895: Pixel = 58;
			7896: Pixel = 76;
			7897: Pixel = 79;
			7898: Pixel = 86;
			7899: Pixel = 86;
			7900: Pixel = 135;
			7901: Pixel = 145;
			7902: Pixel = 128;
			7903: Pixel = 100;
			7904: Pixel = 62;
			7905: Pixel = 55;
			7906: Pixel = 123;
			7907: Pixel = 164;
			7908: Pixel = 171;
			7909: Pixel = 171;
			7910: Pixel = 174;
			7911: Pixel = 151;
			7912: Pixel = 153;
			7913: Pixel = 130;
			7914: Pixel = 61;
			7915: Pixel = 41;
			7916: Pixel = 36;
			7917: Pixel = 68;
			7918: Pixel = 97;
			7919: Pixel = 93;
			7920: Pixel = 91;
			7921: Pixel = 71;
			7922: Pixel = 77;
			7923: Pixel = 75;
			7924: Pixel = 84;
			7925: Pixel = 98;
			7926: Pixel = 64;
			7927: Pixel = 86;
			7928: Pixel = 111;
			7929: Pixel = 134;
			7930: Pixel = 140;
			7931: Pixel = 94;
			7932: Pixel = 89;
			7933: Pixel = 96;
			7934: Pixel = 87;
			7935: Pixel = 45;
			7936: Pixel = 55;
			7937: Pixel = 66;
			7938: Pixel = 52;
			7939: Pixel = 50;
			7940: Pixel = 58;
			7941: Pixel = 58;
			7942: Pixel = 51;
			7943: Pixel = 60;
			7944: Pixel = 75;
			7945: Pixel = 57;
			7946: Pixel = 68;
			7947: Pixel = 106;
			7948: Pixel = 119;
			7949: Pixel = 124;
			7950: Pixel = 125;
			7951: Pixel = 133;
			7952: Pixel = 140;
			7953: Pixel = 142;
			7954: Pixel = 137;
			7955: Pixel = 139;
			7956: Pixel = 149;
			7957: Pixel = 160;
			7958: Pixel = 171;
			7959: Pixel = 182;
			7960: Pixel = 187;
			7961: Pixel = 190;
			7962: Pixel = 194;
			7963: Pixel = 199;
			7964: Pixel = 202;
			7965: Pixel = 218;
			7966: Pixel = 205;
			7967: Pixel = 86;
			7968: Pixel = 56;
			7969: Pixel = 74;
			7970: Pixel = 68;
			7971: Pixel = 73;
			7972: Pixel = 62;
			7973: Pixel = 141;
			7974: Pixel = 145;
			7975: Pixel = 148;
			7976: Pixel = 144;
			7977: Pixel = 142;
			7978: Pixel = 140;
			7979: Pixel = 137;
			7980: Pixel = 132;
			7981: Pixel = 125;
			7982: Pixel = 118;
			7983: Pixel = 107;
			7984: Pixel = 106;
			7985: Pixel = 133;
			7986: Pixel = 92;
			7987: Pixel = 143;
			7988: Pixel = 214;
			7989: Pixel = 209;
			7990: Pixel = 210;
			7991: Pixel = 210;
			7992: Pixel = 152;
			7993: Pixel = 48;
			7994: Pixel = 67;
			7995: Pixel = 88;
			7996: Pixel = 80;
			7997: Pixel = 94;
			7998: Pixel = 92;
			7999: Pixel = 84;
			8000: Pixel = 126;
			8001: Pixel = 146;
			8002: Pixel = 150;
			8003: Pixel = 132;
			8004: Pixel = 77;
			8005: Pixel = 54;
			8006: Pixel = 121;
			8007: Pixel = 165;
			8008: Pixel = 175;
			8009: Pixel = 173;
			8010: Pixel = 175;
			8011: Pixel = 153;
			8012: Pixel = 177;
			8013: Pixel = 119;
			8014: Pixel = 50;
			8015: Pixel = 48;
			8016: Pixel = 51;
			8017: Pixel = 61;
			8018: Pixel = 56;
			8019: Pixel = 71;
			8020: Pixel = 58;
			8021: Pixel = 61;
			8022: Pixel = 71;
			8023: Pixel = 50;
			8024: Pixel = 92;
			8025: Pixel = 66;
			8026: Pixel = 63;
			8027: Pixel = 85;
			8028: Pixel = 96;
			8029: Pixel = 124;
			8030: Pixel = 147;
			8031: Pixel = 101;
			8032: Pixel = 108;
			8033: Pixel = 118;
			8034: Pixel = 97;
			8035: Pixel = 45;
			8036: Pixel = 56;
			8037: Pixel = 66;
			8038: Pixel = 54;
			8039: Pixel = 52;
			8040: Pixel = 60;
			8041: Pixel = 59;
			8042: Pixel = 55;
			8043: Pixel = 66;
			8044: Pixel = 89;
			8045: Pixel = 73;
			8046: Pixel = 57;
			8047: Pixel = 112;
			8048: Pixel = 121;
			8049: Pixel = 118;
			8050: Pixel = 130;
			8051: Pixel = 138;
			8052: Pixel = 138;
			8053: Pixel = 140;
			8054: Pixel = 139;
			8055: Pixel = 144;
			8056: Pixel = 154;
			8057: Pixel = 161;
			8058: Pixel = 166;
			8059: Pixel = 174;
			8060: Pixel = 180;
			8061: Pixel = 185;
			8062: Pixel = 190;
			8063: Pixel = 196;
			8064: Pixel = 203;
			8065: Pixel = 205;
			8066: Pixel = 217;
			8067: Pixel = 210;
			8068: Pixel = 87;
			8069: Pixel = 49;
			8070: Pixel = 65;
			8071: Pixel = 70;
			8072: Pixel = 65;
			8073: Pixel = 146;
			8074: Pixel = 144;
			8075: Pixel = 148;
			8076: Pixel = 144;
			8077: Pixel = 143;
			8078: Pixel = 142;
			8079: Pixel = 139;
			8080: Pixel = 137;
			8081: Pixel = 132;
			8082: Pixel = 128;
			8083: Pixel = 122;
			8084: Pixel = 119;
			8085: Pixel = 130;
			8086: Pixel = 113;
			8087: Pixel = 179;
			8088: Pixel = 215;
			8089: Pixel = 212;
			8090: Pixel = 210;
			8091: Pixel = 194;
			8092: Pixel = 99;
			8093: Pixel = 56;
			8094: Pixel = 96;
			8095: Pixel = 88;
			8096: Pixel = 95;
			8097: Pixel = 109;
			8098: Pixel = 91;
			8099: Pixel = 92;
			8100: Pixel = 81;
			8101: Pixel = 131;
			8102: Pixel = 159;
			8103: Pixel = 158;
			8104: Pixel = 96;
			8105: Pixel = 52;
			8106: Pixel = 123;
			8107: Pixel = 167;
			8108: Pixel = 177;
			8109: Pixel = 176;
			8110: Pixel = 177;
			8111: Pixel = 158;
			8112: Pixel = 155;
			8113: Pixel = 89;
			8114: Pixel = 40;
			8115: Pixel = 43;
			8116: Pixel = 52;
			8117: Pixel = 64;
			8118: Pixel = 55;
			8119: Pixel = 42;
			8120: Pixel = 81;
			8121: Pixel = 67;
			8122: Pixel = 40;
			8123: Pixel = 67;
			8124: Pixel = 58;
			8125: Pixel = 84;
			8126: Pixel = 65;
			8127: Pixel = 75;
			8128: Pixel = 90;
			8129: Pixel = 117;
			8130: Pixel = 124;
			8131: Pixel = 141;
			8132: Pixel = 110;
			8133: Pixel = 100;
			8134: Pixel = 123;
			8135: Pixel = 55;
			8136: Pixel = 46;
			8137: Pixel = 67;
			8138: Pixel = 53;
			8139: Pixel = 46;
			8140: Pixel = 57;
			8141: Pixel = 60;
			8142: Pixel = 49;
			8143: Pixel = 61;
			8144: Pixel = 103;
			8145: Pixel = 93;
			8146: Pixel = 51;
			8147: Pixel = 107;
			8148: Pixel = 119;
			8149: Pixel = 130;
			8150: Pixel = 134;
			8151: Pixel = 138;
			8152: Pixel = 139;
			8153: Pixel = 139;
			8154: Pixel = 141;
			8155: Pixel = 145;
			8156: Pixel = 152;
			8157: Pixel = 159;
			8158: Pixel = 163;
			8159: Pixel = 170;
			8160: Pixel = 175;
			8161: Pixel = 180;
			8162: Pixel = 186;
			8163: Pixel = 194;
			8164: Pixel = 200;
			8165: Pixel = 206;
			8166: Pixel = 207;
			8167: Pixel = 223;
			8168: Pixel = 196;
			8169: Pixel = 54;
			8170: Pixel = 52;
			8171: Pixel = 57;
			8172: Pixel = 71;
			8173: Pixel = 147;
			8174: Pixel = 143;
			8175: Pixel = 148;
			8176: Pixel = 144;
			8177: Pixel = 143;
			8178: Pixel = 142;
			8179: Pixel = 141;
			8180: Pixel = 138;
			8181: Pixel = 135;
			8182: Pixel = 131;
			8183: Pixel = 126;
			8184: Pixel = 128;
			8185: Pixel = 133;
			8186: Pixel = 132;
			8187: Pixel = 200;
			8188: Pixel = 215;
			8189: Pixel = 211;
			8190: Pixel = 210;
			8191: Pixel = 158;
			8192: Pixel = 76;
			8193: Pixel = 89;
			8194: Pixel = 93;
			8195: Pixel = 96;
			8196: Pixel = 112;
			8197: Pixel = 102;
			8198: Pixel = 93;
			8199: Pixel = 101;
			8200: Pixel = 40;
			8201: Pixel = 104;
			8202: Pixel = 166;
			8203: Pixel = 167;
			8204: Pixel = 113;
			8205: Pixel = 45;
			8206: Pixel = 120;
			8207: Pixel = 168;
			8208: Pixel = 176;
			8209: Pixel = 177;
			8210: Pixel = 177;
			8211: Pixel = 157;
			8212: Pixel = 144;
			8213: Pixel = 94;
			8214: Pixel = 39;
			8215: Pixel = 43;
			8216: Pixel = 61;
			8217: Pixel = 54;
			8218: Pixel = 48;
			8219: Pixel = 47;
			8220: Pixel = 93;
			8221: Pixel = 67;
			8222: Pixel = 46;
			8223: Pixel = 56;
			8224: Pixel = 71;
			8225: Pixel = 74;
			8226: Pixel = 80;
			8227: Pixel = 94;
			8228: Pixel = 87;
			8229: Pixel = 95;
			8230: Pixel = 116;
			8231: Pixel = 153;
			8232: Pixel = 106;
			8233: Pixel = 51;
			8234: Pixel = 158;
			8235: Pixel = 71;
			8236: Pixel = 36;
			8237: Pixel = 67;
			8238: Pixel = 55;
			8239: Pixel = 45;
			8240: Pixel = 58;
			8241: Pixel = 60;
			8242: Pixel = 49;
			8243: Pixel = 58;
			8244: Pixel = 111;
			8245: Pixel = 97;
			8246: Pixel = 48;
			8247: Pixel = 102;
			8248: Pixel = 127;
			8249: Pixel = 133;
			8250: Pixel = 132;
			8251: Pixel = 136;
			8252: Pixel = 140;
			8253: Pixel = 140;
			8254: Pixel = 142;
			8255: Pixel = 146;
			8256: Pixel = 150;
			8257: Pixel = 156;
			8258: Pixel = 161;
			8259: Pixel = 166;
			8260: Pixel = 173;
			8261: Pixel = 179;
			8262: Pixel = 184;
			8263: Pixel = 191;
			8264: Pixel = 198;
			8265: Pixel = 204;
			8266: Pixel = 208;
			8267: Pixel = 210;
			8268: Pixel = 233;
			8269: Pixel = 139;
			8270: Pixel = 38;
			8271: Pixel = 45;
			8272: Pixel = 78;
			8273: Pixel = 148;
			8274: Pixel = 143;
			8275: Pixel = 146;
			8276: Pixel = 144;
			8277: Pixel = 143;
			8278: Pixel = 141;
			8279: Pixel = 140;
			8280: Pixel = 138;
			8281: Pixel = 137;
			8282: Pixel = 132;
			8283: Pixel = 126;
			8284: Pixel = 124;
			8285: Pixel = 144;
			8286: Pixel = 168;
			8287: Pixel = 208;
			8288: Pixel = 215;
			8289: Pixel = 211;
			8290: Pixel = 204;
			8291: Pixel = 117;
			8292: Pixel = 79;
			8293: Pixel = 93;
			8294: Pixel = 98;
			8295: Pixel = 110;
			8296: Pixel = 103;
			8297: Pixel = 88;
			8298: Pixel = 101;
			8299: Pixel = 103;
			8300: Pixel = 33;
			8301: Pixel = 85;
			8302: Pixel = 166;
			8303: Pixel = 174;
			8304: Pixel = 114;
			8305: Pixel = 38;
			8306: Pixel = 118;
			8307: Pixel = 168;
			8308: Pixel = 178;
			8309: Pixel = 176;
			8310: Pixel = 179;
			8311: Pixel = 162;
			8312: Pixel = 133;
			8313: Pixel = 96;
			8314: Pixel = 40;
			8315: Pixel = 50;
			8316: Pixel = 56;
			8317: Pixel = 46;
			8318: Pixel = 48;
			8319: Pixel = 50;
			8320: Pixel = 105;
			8321: Pixel = 56;
			8322: Pixel = 57;
			8323: Pixel = 42;
			8324: Pixel = 69;
			8325: Pixel = 66;
			8326: Pixel = 69;
			8327: Pixel = 101;
			8328: Pixel = 99;
			8329: Pixel = 78;
			8330: Pixel = 124;
			8331: Pixel = 152;
			8332: Pixel = 93;
			8333: Pixel = 46;
			8334: Pixel = 167;
			8335: Pixel = 61;
			8336: Pixel = 43;
			8337: Pixel = 73;
			8338: Pixel = 61;
			8339: Pixel = 46;
			8340: Pixel = 58;
			8341: Pixel = 53;
			8342: Pixel = 47;
			8343: Pixel = 71;
			8344: Pixel = 107;
			8345: Pixel = 96;
			8346: Pixel = 55;
			8347: Pixel = 104;
			8348: Pixel = 129;
			8349: Pixel = 128;
			8350: Pixel = 135;
			8351: Pixel = 137;
			8352: Pixel = 138;
			8353: Pixel = 139;
			8354: Pixel = 143;
			8355: Pixel = 146;
			8356: Pixel = 148;
			8357: Pixel = 154;
			8358: Pixel = 158;
			8359: Pixel = 164;
			8360: Pixel = 171;
			8361: Pixel = 176;
			8362: Pixel = 183;
			8363: Pixel = 188;
			8364: Pixel = 197;
			8365: Pixel = 204;
			8366: Pixel = 209;
			8367: Pixel = 212;
			8368: Pixel = 221;
			8369: Pixel = 211;
			8370: Pixel = 60;
			8371: Pixel = 26;
			8372: Pixel = 88;
			8373: Pixel = 152;
			8374: Pixel = 145;
			8375: Pixel = 148;
			8376: Pixel = 145;
			8377: Pixel = 144;
			8378: Pixel = 141;
			8379: Pixel = 137;
			8380: Pixel = 135;
			8381: Pixel = 134;
			8382: Pixel = 128;
			8383: Pixel = 120;
			8384: Pixel = 142;
			8385: Pixel = 186;
			8386: Pixel = 201;
			8387: Pixel = 213;
			8388: Pixel = 214;
			8389: Pixel = 213;
			8390: Pixel = 175;
			8391: Pixel = 94;
			8392: Pixel = 92;
			8393: Pixel = 96;
			8394: Pixel = 108;
			8395: Pixel = 109;
			8396: Pixel = 90;
			8397: Pixel = 94;
			8398: Pixel = 102;
			8399: Pixel = 101;
			8400: Pixel = 29;
			8401: Pixel = 74;
			8402: Pixel = 158;
			8403: Pixel = 174;
			8404: Pixel = 113;
			8405: Pixel = 36;
			8406: Pixel = 116;
			8407: Pixel = 169;
			8408: Pixel = 178;
			8409: Pixel = 178;
			8410: Pixel = 181;
			8411: Pixel = 161;
			8412: Pixel = 148;
			8413: Pixel = 77;
			8414: Pixel = 43;
			8415: Pixel = 55;
			8416: Pixel = 46;
			8417: Pixel = 47;
			8418: Pixel = 37;
			8419: Pixel = 76;
			8420: Pixel = 116;
			8421: Pixel = 41;
			8422: Pixel = 54;
			8423: Pixel = 59;
			8424: Pixel = 49;
			8425: Pixel = 46;
			8426: Pixel = 61;
			8427: Pixel = 88;
			8428: Pixel = 104;
			8429: Pixel = 64;
			8430: Pixel = 119;
			8431: Pixel = 145;
			8432: Pixel = 117;
			8433: Pixel = 71;
			8434: Pixel = 149;
			8435: Pixel = 77;
			8436: Pixel = 50;
			8437: Pixel = 73;
			8438: Pixel = 59;
			8439: Pixel = 50;
			8440: Pixel = 54;
			8441: Pixel = 54;
			8442: Pixel = 51;
			8443: Pixel = 84;
			8444: Pixel = 118;
			8445: Pixel = 109;
			8446: Pixel = 60;
			8447: Pixel = 107;
			8448: Pixel = 131;
			8449: Pixel = 132;
			8450: Pixel = 136;
			8451: Pixel = 137;
			8452: Pixel = 136;
			8453: Pixel = 136;
			8454: Pixel = 140;
			8455: Pixel = 144;
			8456: Pixel = 146;
			8457: Pixel = 152;
			8458: Pixel = 156;
			8459: Pixel = 163;
			8460: Pixel = 167;
			8461: Pixel = 174;
			8462: Pixel = 181;
			8463: Pixel = 188;
			8464: Pixel = 195;
			8465: Pixel = 203;
			8466: Pixel = 209;
			8467: Pixel = 212;
			8468: Pixel = 212;
			8469: Pixel = 232;
			8470: Pixel = 121;
			8471: Pixel = 14;
			8472: Pixel = 100;
			8473: Pixel = 152;
			8474: Pixel = 146;
			8475: Pixel = 146;
			8476: Pixel = 145;
			8477: Pixel = 143;
			8478: Pixel = 140;
			8479: Pixel = 136;
			8480: Pixel = 133;
			8481: Pixel = 130;
			8482: Pixel = 125;
			8483: Pixel = 124;
			8484: Pixel = 189;
			8485: Pixel = 213;
			8486: Pixel = 204;
			8487: Pixel = 215;
			8488: Pixel = 216;
			8489: Pixel = 205;
			8490: Pixel = 133;
			8491: Pixel = 88;
			8492: Pixel = 92;
			8493: Pixel = 104;
			8494: Pixel = 116;
			8495: Pixel = 100;
			8496: Pixel = 89;
			8497: Pixel = 103;
			8498: Pixel = 102;
			8499: Pixel = 101;
			8500: Pixel = 27;
			8501: Pixel = 63;
			8502: Pixel = 155;
			8503: Pixel = 176;
			8504: Pixel = 122;
			8505: Pixel = 38;
			8506: Pixel = 113;
			8507: Pixel = 170;
			8508: Pixel = 178;
			8509: Pixel = 178;
			8510: Pixel = 179;
			8511: Pixel = 164;
			8512: Pixel = 133;
			8513: Pixel = 61;
			8514: Pixel = 54;
			8515: Pixel = 46;
			8516: Pixel = 44;
			8517: Pixel = 44;
			8518: Pixel = 53;
			8519: Pixel = 95;
			8520: Pixel = 89;
			8521: Pixel = 40;
			8522: Pixel = 57;
			8523: Pixel = 58;
			8524: Pixel = 41;
			8525: Pixel = 53;
			8526: Pixel = 53;
			8527: Pixel = 66;
			8528: Pixel = 106;
			8529: Pixel = 85;
			8530: Pixel = 128;
			8531: Pixel = 138;
			8532: Pixel = 122;
			8533: Pixel = 155;
			8534: Pixel = 124;
			8535: Pixel = 68;
			8536: Pixel = 51;
			8537: Pixel = 55;
			8538: Pixel = 56;
			8539: Pixel = 56;
			8540: Pixel = 53;
			8541: Pixel = 51;
			8542: Pixel = 66;
			8543: Pixel = 109;
			8544: Pixel = 130;
			8545: Pixel = 103;
			8546: Pixel = 64;
			8547: Pixel = 111;
			8548: Pixel = 129;
			8549: Pixel = 134;
			8550: Pixel = 138;
			8551: Pixel = 137;
			8552: Pixel = 136;
			8553: Pixel = 137;
			8554: Pixel = 140;
			8555: Pixel = 143;
			8556: Pixel = 145;
			8557: Pixel = 149;
			8558: Pixel = 156;
			8559: Pixel = 160;
			8560: Pixel = 164;
			8561: Pixel = 173;
			8562: Pixel = 179;
			8563: Pixel = 186;
			8564: Pixel = 194;
			8565: Pixel = 201;
			8566: Pixel = 207;
			8567: Pixel = 210;
			8568: Pixel = 211;
			8569: Pixel = 227;
			8570: Pixel = 176;
			8571: Pixel = 21;
			8572: Pixel = 108;
			8573: Pixel = 151;
			8574: Pixel = 147;
			8575: Pixel = 144;
			8576: Pixel = 143;
			8577: Pixel = 141;
			8578: Pixel = 139;
			8579: Pixel = 137;
			8580: Pixel = 133;
			8581: Pixel = 129;
			8582: Pixel = 120;
			8583: Pixel = 135;
			8584: Pixel = 209;
			8585: Pixel = 215;
			8586: Pixel = 209;
			8587: Pixel = 216;
			8588: Pixel = 216;
			8589: Pixel = 179;
			8590: Pixel = 111;
			8591: Pixel = 95;
			8592: Pixel = 93;
			8593: Pixel = 109;
			8594: Pixel = 111;
			8595: Pixel = 93;
			8596: Pixel = 97;
			8597: Pixel = 105;
			8598: Pixel = 100;
			8599: Pixel = 90;
			8600: Pixel = 27;
			8601: Pixel = 60;
			8602: Pixel = 152;
			8603: Pixel = 175;
			8604: Pixel = 131;
			8605: Pixel = 44;
			8606: Pixel = 108;
			8607: Pixel = 170;
			8608: Pixel = 176;
			8609: Pixel = 172;
			8610: Pixel = 174;
			8611: Pixel = 161;
			8612: Pixel = 137;
			8613: Pixel = 78;
			8614: Pixel = 44;
			8615: Pixel = 45;
			8616: Pixel = 47;
			8617: Pixel = 56;
			8618: Pixel = 63;
			8619: Pixel = 55;
			8620: Pixel = 85;
			8621: Pixel = 50;
			8622: Pixel = 58;
			8623: Pixel = 53;
			8624: Pixel = 44;
			8625: Pixel = 54;
			8626: Pixel = 64;
			8627: Pixel = 65;
			8628: Pixel = 50;
			8629: Pixel = 121;
			8630: Pixel = 136;
			8631: Pixel = 116;
			8632: Pixel = 82;
			8633: Pixel = 119;
			8634: Pixel = 110;
			8635: Pixel = 92;
			8636: Pixel = 89;
			8637: Pixel = 79;
			8638: Pixel = 72;
			8639: Pixel = 55;
			8640: Pixel = 53;
			8641: Pixel = 51;
			8642: Pixel = 81;
			8643: Pixel = 119;
			8644: Pixel = 130;
			8645: Pixel = 97;
			8646: Pixel = 68;
			8647: Pixel = 117;
			8648: Pixel = 131;
			8649: Pixel = 132;
			8650: Pixel = 140;
			8651: Pixel = 140;
			8652: Pixel = 136;
			8653: Pixel = 134;
			8654: Pixel = 137;
			8655: Pixel = 140;
			8656: Pixel = 143;
			8657: Pixel = 148;
			8658: Pixel = 153;
			8659: Pixel = 158;
			8660: Pixel = 162;
			8661: Pixel = 168;
			8662: Pixel = 175;
			8663: Pixel = 186;
			8664: Pixel = 192;
			8665: Pixel = 199;
			8666: Pixel = 205;
			8667: Pixel = 208;
			8668: Pixel = 211;
			8669: Pixel = 218;
			8670: Pixel = 212;
			8671: Pixel = 53;
			8672: Pixel = 110;
			8673: Pixel = 150;
			8674: Pixel = 147;
			8675: Pixel = 142;
			8676: Pixel = 142;
			8677: Pixel = 139;
			8678: Pixel = 139;
			8679: Pixel = 138;
			8680: Pixel = 134;
			8681: Pixel = 128;
			8682: Pixel = 120;
			8683: Pixel = 148;
			8684: Pixel = 212;
			8685: Pixel = 207;
			8686: Pixel = 208;
			8687: Pixel = 218;
			8688: Pixel = 206;
			8689: Pixel = 145;
			8690: Pixel = 112;
			8691: Pixel = 101;
			8692: Pixel = 98;
			8693: Pixel = 110;
			8694: Pixel = 104;
			8695: Pixel = 89;
			8696: Pixel = 102;
			8697: Pixel = 102;
			8698: Pixel = 92;
			8699: Pixel = 84;
			8700: Pixel = 29;
			8701: Pixel = 51;
			8702: Pixel = 142;
			8703: Pixel = 177;
			8704: Pixel = 136;
			8705: Pixel = 46;
			8706: Pixel = 107;
			8707: Pixel = 168;
			8708: Pixel = 177;
			8709: Pixel = 177;
			8710: Pixel = 178;
			8711: Pixel = 163;
			8712: Pixel = 140;
			8713: Pixel = 66;
			8714: Pixel = 46;
			8715: Pixel = 47;
			8716: Pixel = 45;
			8717: Pixel = 49;
			8718: Pixel = 55;
			8719: Pixel = 54;
			8720: Pixel = 70;
			8721: Pixel = 55;
			8722: Pixel = 49;
			8723: Pixel = 58;
			8724: Pixel = 44;
			8725: Pixel = 47;
			8726: Pixel = 73;
			8727: Pixel = 65;
			8728: Pixel = 59;
			8729: Pixel = 99;
			8730: Pixel = 117;
			8731: Pixel = 122;
			8732: Pixel = 92;
			8733: Pixel = 49;
			8734: Pixel = 50;
			8735: Pixel = 58;
			8736: Pixel = 75;
			8737: Pixel = 89;
			8738: Pixel = 87;
			8739: Pixel = 59;
			8740: Pixel = 47;
			8741: Pixel = 63;
			8742: Pixel = 97;
			8743: Pixel = 123;
			8744: Pixel = 133;
			8745: Pixel = 91;
			8746: Pixel = 79;
			8747: Pixel = 126;
			8748: Pixel = 133;
			8749: Pixel = 136;
			8750: Pixel = 139;
			8751: Pixel = 140;
			8752: Pixel = 138;
			8753: Pixel = 134;
			8754: Pixel = 136;
			8755: Pixel = 139;
			8756: Pixel = 142;
			8757: Pixel = 147;
			8758: Pixel = 151;
			8759: Pixel = 156;
			8760: Pixel = 160;
			8761: Pixel = 167;
			8762: Pixel = 172;
			8763: Pixel = 182;
			8764: Pixel = 191;
			8765: Pixel = 197;
			8766: Pixel = 203;
			8767: Pixel = 207;
			8768: Pixel = 210;
			8769: Pixel = 212;
			8770: Pixel = 225;
			8771: Pixel = 101;
			8772: Pixel = 111;
			8773: Pixel = 151;
			8774: Pixel = 147;
			8775: Pixel = 142;
			8776: Pixel = 142;
			8777: Pixel = 138;
			8778: Pixel = 139;
			8779: Pixel = 138;
			8780: Pixel = 134;
			8781: Pixel = 128;
			8782: Pixel = 124;
			8783: Pixel = 150;
			8784: Pixel = 211;
			8785: Pixel = 206;
			8786: Pixel = 209;
			8787: Pixel = 219;
			8788: Pixel = 185;
			8789: Pixel = 123;
			8790: Pixel = 113;
			8791: Pixel = 100;
			8792: Pixel = 97;
			8793: Pixel = 104;
			8794: Pixel = 88;
			8795: Pixel = 93;
			8796: Pixel = 104;
			8797: Pixel = 96;
			8798: Pixel = 91;
			8799: Pixel = 93;
			8800: Pixel = 35;
			8801: Pixel = 44;
			8802: Pixel = 131;
			8803: Pixel = 175;
			8804: Pixel = 141;
			8805: Pixel = 57;
			8806: Pixel = 105;
			8807: Pixel = 166;
			8808: Pixel = 177;
			8809: Pixel = 177;
			8810: Pixel = 178;
			8811: Pixel = 161;
			8812: Pixel = 147;
			8813: Pixel = 76;
			8814: Pixel = 48;
			8815: Pixel = 41;
			8816: Pixel = 55;
			8817: Pixel = 69;
			8818: Pixel = 53;
			8819: Pixel = 50;
			8820: Pixel = 61;
			8821: Pixel = 53;
			8822: Pixel = 51;
			8823: Pixel = 59;
			8824: Pixel = 49;
			8825: Pixel = 54;
			8826: Pixel = 69;
			8827: Pixel = 74;
			8828: Pixel = 74;
			8829: Pixel = 110;
			8830: Pixel = 124;
			8831: Pixel = 87;
			8832: Pixel = 114;
			8833: Pixel = 106;
			8834: Pixel = 66;
			8835: Pixel = 48;
			8836: Pixel = 52;
			8837: Pixel = 52;
			8838: Pixel = 54;
			8839: Pixel = 53;
			8840: Pixel = 46;
			8841: Pixel = 77;
			8842: Pixel = 107;
			8843: Pixel = 123;
			8844: Pixel = 128;
			8845: Pixel = 76;
			8846: Pixel = 92;
			8847: Pixel = 131;
			8848: Pixel = 137;
			8849: Pixel = 140;
			8850: Pixel = 141;
			8851: Pixel = 140;
			8852: Pixel = 138;
			8853: Pixel = 135;
			8854: Pixel = 136;
			8855: Pixel = 137;
			8856: Pixel = 141;
			8857: Pixel = 146;
			8858: Pixel = 149;
			8859: Pixel = 154;
			8860: Pixel = 159;
			8861: Pixel = 164;
			8862: Pixel = 168;
			8863: Pixel = 178;
			8864: Pixel = 188;
			8865: Pixel = 195;
			8866: Pixel = 200;
			8867: Pixel = 206;
			8868: Pixel = 209;
			8869: Pixel = 210;
			8870: Pixel = 223;
			8871: Pixel = 156;
			8872: Pixel = 120;
			8873: Pixel = 146;
			8874: Pixel = 144;
			8875: Pixel = 143;
			8876: Pixel = 145;
			8877: Pixel = 144;
			8878: Pixel = 141;
			8879: Pixel = 140;
			8880: Pixel = 134;
			8881: Pixel = 131;
			8882: Pixel = 134;
			8883: Pixel = 138;
			8884: Pixel = 168;
			8885: Pixel = 187;
			8886: Pixel = 212;
			8887: Pixel = 216;
			8888: Pixel = 169;
			8889: Pixel = 113;
			8890: Pixel = 108;
			8891: Pixel = 95;
			8892: Pixel = 99;
			8893: Pixel = 85;
			8894: Pixel = 85;
			8895: Pixel = 107;
			8896: Pixel = 95;
			8897: Pixel = 91;
			8898: Pixel = 95;
			8899: Pixel = 94;
			8900: Pixel = 37;
			8901: Pixel = 39;
			8902: Pixel = 122;
			8903: Pixel = 170;
			8904: Pixel = 145;
			8905: Pixel = 68;
			8906: Pixel = 103;
			8907: Pixel = 164;
			8908: Pixel = 175;
			8909: Pixel = 175;
			8910: Pixel = 178;
			8911: Pixel = 161;
			8912: Pixel = 145;
			8913: Pixel = 91;
			8914: Pixel = 50;
			8915: Pixel = 44;
			8916: Pixel = 64;
			8917: Pixel = 53;
			8918: Pixel = 43;
			8919: Pixel = 58;
			8920: Pixel = 61;
			8921: Pixel = 59;
			8922: Pixel = 60;
			8923: Pixel = 56;
			8924: Pixel = 50;
			8925: Pixel = 66;
			8926: Pixel = 53;
			8927: Pixel = 72;
			8928: Pixel = 77;
			8929: Pixel = 63;
			8930: Pixel = 99;
			8931: Pixel = 89;
			8932: Pixel = 63;
			8933: Pixel = 145;
			8934: Pixel = 101;
			8935: Pixel = 42;
			8936: Pixel = 52;
			8937: Pixel = 54;
			8938: Pixel = 47;
			8939: Pixel = 44;
			8940: Pixel = 55;
			8941: Pixel = 90;
			8942: Pixel = 115;
			8943: Pixel = 126;
			8944: Pixel = 114;
			8945: Pixel = 66;
			8946: Pixel = 111;
			8947: Pixel = 135;
			8948: Pixel = 138;
			8949: Pixel = 139;
			8950: Pixel = 143;
			8951: Pixel = 141;
			8952: Pixel = 139;
			8953: Pixel = 138;
			8954: Pixel = 135;
			8955: Pixel = 138;
			8956: Pixel = 141;
			8957: Pixel = 145;
			8958: Pixel = 149;
			8959: Pixel = 151;
			8960: Pixel = 155;
			8961: Pixel = 160;
			8962: Pixel = 167;
			8963: Pixel = 175;
			8964: Pixel = 184;
			8965: Pixel = 192;
			8966: Pixel = 199;
			8967: Pixel = 205;
			8968: Pixel = 210;
			8969: Pixel = 211;
			8970: Pixel = 216;
			8971: Pixel = 200;
			8972: Pixel = 136;
			8973: Pixel = 107;
			8974: Pixel = 112;
			8975: Pixel = 125;
			8976: Pixel = 137;
			8977: Pixel = 143;
			8978: Pixel = 145;
			8979: Pixel = 143;
			8980: Pixel = 139;
			8981: Pixel = 137;
			8982: Pixel = 145;
			8983: Pixel = 144;
			8984: Pixel = 130;
			8985: Pixel = 168;
			8986: Pixel = 219;
			8987: Pixel = 210;
			8988: Pixel = 151;
			8989: Pixel = 108;
			8990: Pixel = 96;
			8991: Pixel = 94;
			8992: Pixel = 93;
			8993: Pixel = 78;
			8994: Pixel = 100;
			8995: Pixel = 101;
			8996: Pixel = 88;
			8997: Pixel = 93;
			8998: Pixel = 96;
			8999: Pixel = 81;
			9000: Pixel = 34;
			9001: Pixel = 37;
			9002: Pixel = 116;
			9003: Pixel = 175;
			9004: Pixel = 153;
			9005: Pixel = 71;
			9006: Pixel = 99;
			9007: Pixel = 161;
			9008: Pixel = 173;
			9009: Pixel = 176;
			9010: Pixel = 178;
			9011: Pixel = 165;
			9012: Pixel = 134;
			9013: Pixel = 90;
			9014: Pixel = 53;
			9015: Pixel = 46;
			9016: Pixel = 50;
			9017: Pixel = 44;
			9018: Pixel = 54;
			9019: Pixel = 61;
			9020: Pixel = 54;
			9021: Pixel = 68;
			9022: Pixel = 52;
			9023: Pixel = 46;
			9024: Pixel = 43;
			9025: Pixel = 55;
			9026: Pixel = 59;
			9027: Pixel = 92;
			9028: Pixel = 120;
			9029: Pixel = 54;
			9030: Pixel = 50;
			9031: Pixel = 68;
			9032: Pixel = 81;
			9033: Pixel = 104;
			9034: Pixel = 58;
			9035: Pixel = 45;
			9036: Pixel = 47;
			9037: Pixel = 48;
			9038: Pixel = 40;
			9039: Pixel = 50;
			9040: Pixel = 71;
			9041: Pixel = 105;
			9042: Pixel = 117;
			9043: Pixel = 128;
			9044: Pixel = 85;
			9045: Pixel = 71;
			9046: Pixel = 129;
			9047: Pixel = 135;
			9048: Pixel = 137;
			9049: Pixel = 141;
			9050: Pixel = 143;
			9051: Pixel = 141;
			9052: Pixel = 142;
			9053: Pixel = 139;
			9054: Pixel = 136;
			9055: Pixel = 137;
			9056: Pixel = 139;
			9057: Pixel = 144;
			9058: Pixel = 147;
			9059: Pixel = 151;
			9060: Pixel = 154;
			9061: Pixel = 160;
			9062: Pixel = 166;
			9063: Pixel = 170;
			9064: Pixel = 180;
			9065: Pixel = 189;
			9066: Pixel = 196;
			9067: Pixel = 204;
			9068: Pixel = 209;
			9069: Pixel = 212;
			9070: Pixel = 213;
			9071: Pixel = 221;
			9072: Pixel = 126;
			9073: Pixel = 70;
			9074: Pixel = 78;
			9075: Pixel = 84;
			9076: Pixel = 97;
			9077: Pixel = 109;
			9078: Pixel = 120;
			9079: Pixel = 128;
			9080: Pixel = 136;
			9081: Pixel = 149;
			9082: Pixel = 157;
			9083: Pixel = 135;
			9084: Pixel = 132;
			9085: Pixel = 188;
			9086: Pixel = 222;
			9087: Pixel = 194;
			9088: Pixel = 129;
			9089: Pixel = 92;
			9090: Pixel = 83;
			9091: Pixel = 96;
			9092: Pixel = 75;
			9093: Pixel = 91;
			9094: Pixel = 101;
			9095: Pixel = 92;
			9096: Pixel = 93;
			9097: Pixel = 102;
			9098: Pixel = 87;
			9099: Pixel = 62;
			9100: Pixel = 34;
			9101: Pixel = 29;
			9102: Pixel = 109;
			9103: Pixel = 179;
			9104: Pixel = 165;
			9105: Pixel = 83;
			9106: Pixel = 93;
			9107: Pixel = 160;
			9108: Pixel = 173;
			9109: Pixel = 175;
			9110: Pixel = 178;
			9111: Pixel = 169;
			9112: Pixel = 123;
			9113: Pixel = 94;
			9114: Pixel = 56;
			9115: Pixel = 46;
			9116: Pixel = 43;
			9117: Pixel = 51;
			9118: Pixel = 59;
			9119: Pixel = 56;
			9120: Pixel = 52;
			9121: Pixel = 62;
			9122: Pixel = 61;
			9123: Pixel = 46;
			9124: Pixel = 49;
			9125: Pixel = 53;
			9126: Pixel = 52;
			9127: Pixel = 77;
			9128: Pixel = 126;
			9129: Pixel = 117;
			9130: Pixel = 76;
			9131: Pixel = 91;
			9132: Pixel = 76;
			9133: Pixel = 53;
			9134: Pixel = 53;
			9135: Pixel = 45;
			9136: Pixel = 45;
			9137: Pixel = 43;
			9138: Pixel = 42;
			9139: Pixel = 59;
			9140: Pixel = 90;
			9141: Pixel = 116;
			9142: Pixel = 121;
			9143: Pixel = 108;
			9144: Pixel = 50;
			9145: Pixel = 103;
			9146: Pixel = 135;
			9147: Pixel = 134;
			9148: Pixel = 137;
			9149: Pixel = 141;
			9150: Pixel = 142;
			9151: Pixel = 141;
			9152: Pixel = 141;
			9153: Pixel = 139;
			9154: Pixel = 137;
			9155: Pixel = 134;
			9156: Pixel = 137;
			9157: Pixel = 141;
			9158: Pixel = 144;
			9159: Pixel = 148;
			9160: Pixel = 152;
			9161: Pixel = 157;
			9162: Pixel = 163;
			9163: Pixel = 168;
			9164: Pixel = 175;
			9165: Pixel = 186;
			9166: Pixel = 194;
			9167: Pixel = 202;
			9168: Pixel = 207;
			9169: Pixel = 211;
			9170: Pixel = 211;
			9171: Pixel = 227;
			9172: Pixel = 143;
			9173: Pixel = 76;
			9174: Pixel = 90;
			9175: Pixel = 81;
			9176: Pixel = 76;
			9177: Pixel = 70;
			9178: Pixel = 70;
			9179: Pixel = 74;
			9180: Pixel = 87;
			9181: Pixel = 121;
			9182: Pixel = 147;
			9183: Pixel = 161;
			9184: Pixel = 153;
			9185: Pixel = 204;
			9186: Pixel = 218;
			9187: Pixel = 163;
			9188: Pixel = 93;
			9189: Pixel = 66;
			9190: Pixel = 83;
			9191: Pixel = 82;
			9192: Pixel = 86;
			9193: Pixel = 103;
			9194: Pixel = 92;
			9195: Pixel = 91;
			9196: Pixel = 98;
			9197: Pixel = 100;
			9198: Pixel = 77;
			9199: Pixel = 53;
			9200: Pixel = 56;
			9201: Pixel = 54;
			9202: Pixel = 107;
			9203: Pixel = 178;
			9204: Pixel = 176;
			9205: Pixel = 93;
			9206: Pixel = 94;
			9207: Pixel = 159;
			9208: Pixel = 174;
			9209: Pixel = 174;
			9210: Pixel = 180;
			9211: Pixel = 168;
			9212: Pixel = 114;
			9213: Pixel = 89;
			9214: Pixel = 48;
			9215: Pixel = 47;
			9216: Pixel = 49;
			9217: Pixel = 55;
			9218: Pixel = 53;
			9219: Pixel = 52;
			9220: Pixel = 55;
			9221: Pixel = 63;
			9222: Pixel = 59;
			9223: Pixel = 55;
			9224: Pixel = 46;
			9225: Pixel = 49;
			9226: Pixel = 51;
			9227: Pixel = 45;
			9228: Pixel = 82;
			9229: Pixel = 143;
			9230: Pixel = 122;
			9231: Pixel = 99;
			9232: Pixel = 81;
			9233: Pixel = 40;
			9234: Pixel = 49;
			9235: Pixel = 45;
			9236: Pixel = 43;
			9237: Pixel = 39;
			9238: Pixel = 46;
			9239: Pixel = 75;
			9240: Pixel = 104;
			9241: Pixel = 117;
			9242: Pixel = 122;
			9243: Pixel = 57;
			9244: Pixel = 70;
			9245: Pixel = 130;
			9246: Pixel = 135;
			9247: Pixel = 136;
			9248: Pixel = 138;
			9249: Pixel = 138;
			9250: Pixel = 140;
			9251: Pixel = 143;
			9252: Pixel = 143;
			9253: Pixel = 141;
			9254: Pixel = 139;
			9255: Pixel = 136;
			9256: Pixel = 137;
			9257: Pixel = 138;
			9258: Pixel = 141;
			9259: Pixel = 146;
			9260: Pixel = 151;
			9261: Pixel = 155;
			9262: Pixel = 158;
			9263: Pixel = 165;
			9264: Pixel = 175;
			9265: Pixel = 182;
			9266: Pixel = 191;
			9267: Pixel = 199;
			9268: Pixel = 205;
			9269: Pixel = 209;
			9270: Pixel = 211;
			9271: Pixel = 222;
			9272: Pixel = 183;
			9273: Pixel = 86;
			9274: Pixel = 105;
			9275: Pixel = 100;
			9276: Pixel = 91;
			9277: Pixel = 78;
			9278: Pixel = 62;
			9279: Pixel = 46;
			9280: Pixel = 38;
			9281: Pixel = 60;
			9282: Pixel = 168;
			9283: Pixel = 192;
			9284: Pixel = 166;
			9285: Pixel = 213;
			9286: Pixel = 206;
			9287: Pixel = 118;
			9288: Pixel = 60;
			9289: Pixel = 70;
			9290: Pixel = 78;
			9291: Pixel = 79;
			9292: Pixel = 107;
			9293: Pixel = 95;
			9294: Pixel = 84;
			9295: Pixel = 89;
			9296: Pixel = 104;
			9297: Pixel = 93;
			9298: Pixel = 65;
			9299: Pixel = 52;
			9300: Pixel = 90;
			9301: Pixel = 87;
			9302: Pixel = 117;
			9303: Pixel = 174;
			9304: Pixel = 183;
			9305: Pixel = 109;
			9306: Pixel = 96;
			9307: Pixel = 157;
			9308: Pixel = 175;
			9309: Pixel = 176;
			9310: Pixel = 183;
			9311: Pixel = 165;
			9312: Pixel = 117;
			9313: Pixel = 92;
			9314: Pixel = 43;
			9315: Pixel = 52;
			9316: Pixel = 55;
			9317: Pixel = 45;
			9318: Pixel = 51;
			9319: Pixel = 50;
			9320: Pixel = 54;
			9321: Pixel = 59;
			9322: Pixel = 62;
			9323: Pixel = 52;
			9324: Pixel = 45;
			9325: Pixel = 47;
			9326: Pixel = 57;
			9327: Pixel = 59;
			9328: Pixel = 46;
			9329: Pixel = 91;
			9330: Pixel = 129;
			9331: Pixel = 114;
			9332: Pixel = 91;
			9333: Pixel = 46;
			9334: Pixel = 44;
			9335: Pixel = 42;
			9336: Pixel = 39;
			9337: Pixel = 42;
			9338: Pixel = 62;
			9339: Pixel = 91;
			9340: Pixel = 120;
			9341: Pixel = 122;
			9342: Pixel = 65;
			9343: Pixel = 55;
			9344: Pixel = 117;
			9345: Pixel = 133;
			9346: Pixel = 134;
			9347: Pixel = 137;
			9348: Pixel = 138;
			9349: Pixel = 139;
			9350: Pixel = 140;
			9351: Pixel = 142;
			9352: Pixel = 142;
			9353: Pixel = 142;
			9354: Pixel = 139;
			9355: Pixel = 138;
			9356: Pixel = 136;
			9357: Pixel = 139;
			9358: Pixel = 139;
			9359: Pixel = 143;
			9360: Pixel = 147;
			9361: Pixel = 153;
			9362: Pixel = 156;
			9363: Pixel = 163;
			9364: Pixel = 169;
			9365: Pixel = 178;
			9366: Pixel = 189;
			9367: Pixel = 196;
			9368: Pixel = 203;
			9369: Pixel = 207;
			9370: Pixel = 210;
			9371: Pixel = 214;
			9372: Pixel = 210;
			9373: Pixel = 101;
			9374: Pixel = 98;
			9375: Pixel = 109;
			9376: Pixel = 101;
			9377: Pixel = 92;
			9378: Pixel = 80;
			9379: Pixel = 63;
			9380: Pixel = 40;
			9381: Pixel = 56;
			9382: Pixel = 186;
			9383: Pixel = 188;
			9384: Pixel = 180;
			9385: Pixel = 213;
			9386: Pixel = 146;
			9387: Pixel = 56;
			9388: Pixel = 61;
			9389: Pixel = 73;
			9390: Pixel = 73;
			9391: Pixel = 100;
			9392: Pixel = 99;
			9393: Pixel = 78;
			9394: Pixel = 79;
			9395: Pixel = 98;
			9396: Pixel = 110;
			9397: Pixel = 88;
			9398: Pixel = 70;
			9399: Pixel = 59;
			9400: Pixel = 87;
			9401: Pixel = 105;
			9402: Pixel = 131;
			9403: Pixel = 172;
			9404: Pixel = 181;
			9405: Pixel = 120;
			9406: Pixel = 98;
			9407: Pixel = 156;
			9408: Pixel = 175;
			9409: Pixel = 177;
			9410: Pixel = 184;
			9411: Pixel = 164;
			9412: Pixel = 114;
			9413: Pixel = 85;
			9414: Pixel = 44;
			9415: Pixel = 49;
			9416: Pixel = 48;
			9417: Pixel = 49;
			9418: Pixel = 54;
			9419: Pixel = 49;
			9420: Pixel = 47;
			9421: Pixel = 66;
			9422: Pixel = 58;
			9423: Pixel = 71;
			9424: Pixel = 43;
			9425: Pixel = 60;
			9426: Pixel = 66;
			9427: Pixel = 61;
			9428: Pixel = 65;
			9429: Pixel = 73;
			9430: Pixel = 97;
			9431: Pixel = 99;
			9432: Pixel = 67;
			9433: Pixel = 42;
			9434: Pixel = 47;
			9435: Pixel = 40;
			9436: Pixel = 38;
			9437: Pixel = 58;
			9438: Pixel = 86;
			9439: Pixel = 106;
			9440: Pixel = 101;
			9441: Pixel = 58;
			9442: Pixel = 57;
			9443: Pixel = 108;
			9444: Pixel = 128;
			9445: Pixel = 130;
			9446: Pixel = 135;
			9447: Pixel = 138;
			9448: Pixel = 139;
			9449: Pixel = 139;
			9450: Pixel = 139;
			9451: Pixel = 142;
			9452: Pixel = 142;
			9453: Pixel = 143;
			9454: Pixel = 142;
			9455: Pixel = 140;
			9456: Pixel = 138;
			9457: Pixel = 140;
			9458: Pixel = 138;
			9459: Pixel = 142;
			9460: Pixel = 146;
			9461: Pixel = 148;
			9462: Pixel = 155;
			9463: Pixel = 161;
			9464: Pixel = 165;
			9465: Pixel = 172;
			9466: Pixel = 182;
			9467: Pixel = 192;
			9468: Pixel = 199;
			9469: Pixel = 206;
			9470: Pixel = 210;
			9471: Pixel = 210;
			9472: Pixel = 222;
			9473: Pixel = 130;
			9474: Pixel = 85;
			9475: Pixel = 109;
			9476: Pixel = 103;
			9477: Pixel = 96;
			9478: Pixel = 91;
			9479: Pixel = 79;
			9480: Pixel = 68;
			9481: Pixel = 76;
			9482: Pixel = 171;
			9483: Pixel = 213;
			9484: Pixel = 186;
			9485: Pixel = 134;
			9486: Pixel = 65;
			9487: Pixel = 54;
			9488: Pixel = 70;
			9489: Pixel = 68;
			9490: Pixel = 94;
			9491: Pixel = 104;
			9492: Pixel = 80;
			9493: Pixel = 74;
			9494: Pixel = 89;
			9495: Pixel = 111;
			9496: Pixel = 101;
			9497: Pixel = 84;
			9498: Pixel = 66;
			9499: Pixel = 66;
			9500: Pixel = 70;
			9501: Pixel = 103;
			9502: Pixel = 116;
			9503: Pixel = 165;
			9504: Pixel = 179;
			9505: Pixel = 123;
			9506: Pixel = 99;
			9507: Pixel = 154;
			9508: Pixel = 175;
			9509: Pixel = 178;
			9510: Pixel = 183;
			9511: Pixel = 167;
			9512: Pixel = 109;
			9513: Pixel = 71;
			9514: Pixel = 40;
			9515: Pixel = 52;
			9516: Pixel = 55;
			9517: Pixel = 52;
			9518: Pixel = 56;
			9519: Pixel = 52;
			9520: Pixel = 50;
			9521: Pixel = 82;
			9522: Pixel = 61;
			9523: Pixel = 91;
			9524: Pixel = 60;
			9525: Pixel = 57;
			9526: Pixel = 63;
			9527: Pixel = 67;
			9528: Pixel = 74;
			9529: Pixel = 67;
			9530: Pixel = 124;
			9531: Pixel = 85;
			9532: Pixel = 55;
			9533: Pixel = 42;
			9534: Pixel = 45;
			9535: Pixel = 42;
			9536: Pixel = 43;
			9537: Pixel = 62;
			9538: Pixel = 69;
			9539: Pixel = 61;
			9540: Pixel = 57;
			9541: Pixel = 82;
			9542: Pixel = 116;
			9543: Pixel = 122;
			9544: Pixel = 127;
			9545: Pixel = 131;
			9546: Pixel = 135;
			9547: Pixel = 136;
			9548: Pixel = 138;
			9549: Pixel = 140;
			9550: Pixel = 139;
			9551: Pixel = 142;
			9552: Pixel = 143;
			9553: Pixel = 145;
			9554: Pixel = 145;
			9555: Pixel = 143;
			9556: Pixel = 141;
			9557: Pixel = 139;
			9558: Pixel = 139;
			9559: Pixel = 140;
			9560: Pixel = 144;
			9561: Pixel = 148;
			9562: Pixel = 153;
			9563: Pixel = 158;
			9564: Pixel = 164;
			9565: Pixel = 171;
			9566: Pixel = 178;
			9567: Pixel = 187;
			9568: Pixel = 195;
			9569: Pixel = 203;
			9570: Pixel = 209;
			9571: Pixel = 210;
			9572: Pixel = 222;
			9573: Pixel = 164;
			9574: Pixel = 80;
			9575: Pixel = 101;
			9576: Pixel = 103;
			9577: Pixel = 101;
			9578: Pixel = 99;
			9579: Pixel = 92;
			9580: Pixel = 97;
			9581: Pixel = 94;
			9582: Pixel = 166;
			9583: Pixel = 195;
			9584: Pixel = 116;
			9585: Pixel = 69;
			9586: Pixel = 65;
			9587: Pixel = 75;
			9588: Pixel = 72;
			9589: Pixel = 94;
			9590: Pixel = 108;
			9591: Pixel = 86;
			9592: Pixel = 67;
			9593: Pixel = 77;
			9594: Pixel = 106;
			9595: Pixel = 111;
			9596: Pixel = 97;
			9597: Pixel = 71;
			9598: Pixel = 66;
			9599: Pixel = 65;
			9600: Pixel = 52;
			9601: Pixel = 77;
			9602: Pixel = 102;
			9603: Pixel = 156;
			9604: Pixel = 176;
			9605: Pixel = 131;
			9606: Pixel = 102;
			9607: Pixel = 150;
			9608: Pixel = 175;
			9609: Pixel = 180;
			9610: Pixel = 182;
			9611: Pixel = 175;
			9612: Pixel = 103;
			9613: Pixel = 50;
			9614: Pixel = 46;
			9615: Pixel = 49;
			9616: Pixel = 55;
			9617: Pixel = 57;
			9618: Pixel = 63;
			9619: Pixel = 58;
			9620: Pixel = 50;
			9621: Pixel = 76;
			9622: Pixel = 51;
			9623: Pixel = 100;
			9624: Pixel = 93;
			9625: Pixel = 46;
			9626: Pixel = 84;
			9627: Pixel = 50;
			9628: Pixel = 87;
			9629: Pixel = 68;
			9630: Pixel = 115;
			9631: Pixel = 112;
			9632: Pixel = 60;
			9633: Pixel = 44;
			9634: Pixel = 46;
			9635: Pixel = 43;
			9636: Pixel = 46;
			9637: Pixel = 55;
			9638: Pixel = 68;
			9639: Pixel = 85;
			9640: Pixel = 110;
			9641: Pixel = 122;
			9642: Pixel = 124;
			9643: Pixel = 127;
			9644: Pixel = 127;
			9645: Pixel = 128;
			9646: Pixel = 132;
			9647: Pixel = 135;
			9648: Pixel = 137;
			9649: Pixel = 137;
			9650: Pixel = 140;
			9651: Pixel = 141;
			9652: Pixel = 142;
			9653: Pixel = 145;
			9654: Pixel = 146;
			9655: Pixel = 143;
			9656: Pixel = 143;
			9657: Pixel = 141;
			9658: Pixel = 141;
			9659: Pixel = 141;
			9660: Pixel = 142;
			9661: Pixel = 147;
			9662: Pixel = 151;
			9663: Pixel = 157;
			9664: Pixel = 161;
			9665: Pixel = 169;
			9666: Pixel = 178;
			9667: Pixel = 185;
			9668: Pixel = 192;
			9669: Pixel = 199;
			9670: Pixel = 206;
			9671: Pixel = 210;
			9672: Pixel = 217;
			9673: Pixel = 196;
			9674: Pixel = 85;
			9675: Pixel = 91;
			9676: Pixel = 101;
			9677: Pixel = 108;
			9678: Pixel = 104;
			9679: Pixel = 106;
			9680: Pixel = 114;
			9681: Pixel = 108;
			9682: Pixel = 120;
			9683: Pixel = 111;
			9684: Pixel = 80;
			9685: Pixel = 86;
			9686: Pixel = 87;
			9687: Pixel = 74;
			9688: Pixel = 85;
			9689: Pixel = 107;
			9690: Pixel = 89;
			9691: Pixel = 69;
			9692: Pixel = 65;
			9693: Pixel = 96;
			9694: Pixel = 116;
			9695: Pixel = 112;
			9696: Pixel = 89;
			9697: Pixel = 64;
			9698: Pixel = 62;
			9699: Pixel = 54;
			9700: Pixel = 55;
			9701: Pixel = 61;
			9702: Pixel = 83;
			9703: Pixel = 159;
			9704: Pixel = 196;
			9705: Pixel = 152;
			9706: Pixel = 107;
			9707: Pixel = 150;
			9708: Pixel = 176;
			9709: Pixel = 180;
			9710: Pixel = 185;
			9711: Pixel = 165;
			9712: Pixel = 79;
			9713: Pixel = 54;
			9714: Pixel = 50;
			9715: Pixel = 46;
			9716: Pixel = 55;
			9717: Pixel = 58;
			9718: Pixel = 60;
			9719: Pixel = 65;
			9720: Pixel = 47;
			9721: Pixel = 81;
			9722: Pixel = 43;
			9723: Pixel = 84;
			9724: Pixel = 109;
			9725: Pixel = 52;
			9726: Pixel = 96;
			9727: Pixel = 60;
			9728: Pixel = 64;
			9729: Pixel = 82;
			9730: Pixel = 82;
			9731: Pixel = 99;
			9732: Pixel = 54;
			9733: Pixel = 42;
			9734: Pixel = 47;
			9735: Pixel = 45;
			9736: Pixel = 66;
			9737: Pixel = 93;
			9738: Pixel = 111;
			9739: Pixel = 115;
			9740: Pixel = 119;
			9741: Pixel = 124;
			9742: Pixel = 126;
			9743: Pixel = 128;
			9744: Pixel = 128;
			9745: Pixel = 128;
			9746: Pixel = 133;
			9747: Pixel = 135;
			9748: Pixel = 135;
			9749: Pixel = 138;
			9750: Pixel = 139;
			9751: Pixel = 141;
			9752: Pixel = 141;
			9753: Pixel = 144;
			9754: Pixel = 145;
			9755: Pixel = 146;
			9756: Pixel = 145;
			9757: Pixel = 146;
			9758: Pixel = 143;
			9759: Pixel = 143;
			9760: Pixel = 145;
			9761: Pixel = 147;
			9762: Pixel = 149;
			9763: Pixel = 154;
			9764: Pixel = 160;
			9765: Pixel = 166;
			9766: Pixel = 173;
			9767: Pixel = 181;
			9768: Pixel = 187;
			9769: Pixel = 195;
			9770: Pixel = 202;
			9771: Pixel = 208;
			9772: Pixel = 210;
			9773: Pixel = 214;
			9774: Pixel = 102;
			9775: Pixel = 82;
			9776: Pixel = 102;
			9777: Pixel = 109;
			9778: Pixel = 113;
			9779: Pixel = 118;
			9780: Pixel = 117;
			9781: Pixel = 114;
			9782: Pixel = 106;
			9783: Pixel = 97;
			9784: Pixel = 102;
			9785: Pixel = 107;
			9786: Pixel = 88;
			9787: Pixel = 84;
			9788: Pixel = 98;
			9789: Pixel = 82;
			9790: Pixel = 72;
			9791: Pixel = 71;
			9792: Pixel = 82;
			9793: Pixel = 116;
			9794: Pixel = 119;
			9795: Pixel = 102;
			9796: Pixel = 74;
			9797: Pixel = 59;
			9798: Pixel = 54;
			9799: Pixel = 51;
			9800: Pixel = 52;
			9801: Pixel = 52;
			9802: Pixel = 73;
			9803: Pixel = 178;
			9804: Pixel = 209;
			9805: Pixel = 183;
			9806: Pixel = 117;
			9807: Pixel = 148;
			9808: Pixel = 176;
			9809: Pixel = 178;
			9810: Pixel = 183;
			9811: Pixel = 163;
			9812: Pixel = 86;
			9813: Pixel = 48;
			9814: Pixel = 51;
			9815: Pixel = 51;
			9816: Pixel = 57;
			9817: Pixel = 60;
			9818: Pixel = 65;
			9819: Pixel = 62;
			9820: Pixel = 62;
			9821: Pixel = 90;
			9822: Pixel = 49;
			9823: Pixel = 88;
			9824: Pixel = 99;
			9825: Pixel = 90;
			9826: Pixel = 57;
			9827: Pixel = 84;
			9828: Pixel = 52;
			9829: Pixel = 86;
			9830: Pixel = 60;
			9831: Pixel = 93;
			9832: Pixel = 87;
			9833: Pixel = 42;
			9834: Pixel = 42;
			9835: Pixel = 66;
			9836: Pixel = 91;
			9837: Pixel = 107;
			9838: Pixel = 114;
			9839: Pixel = 118;
			9840: Pixel = 119;
			9841: Pixel = 126;
			9842: Pixel = 126;
			9843: Pixel = 126;
			9844: Pixel = 130;
			9845: Pixel = 131;
			9846: Pixel = 130;
			9847: Pixel = 134;
			9848: Pixel = 136;
			9849: Pixel = 136;
			9850: Pixel = 139;
			9851: Pixel = 139;
			9852: Pixel = 140;
			9853: Pixel = 143;
			9854: Pixel = 145;
			9855: Pixel = 146;
			9856: Pixel = 146;
			9857: Pixel = 147;
			9858: Pixel = 147;
			9859: Pixel = 147;
			9860: Pixel = 146;
			9861: Pixel = 149;
			9862: Pixel = 152;
			9863: Pixel = 153;
			9864: Pixel = 161;
			9865: Pixel = 165;
			9866: Pixel = 171;
			9867: Pixel = 178;
			9868: Pixel = 185;
			9869: Pixel = 193;
			9870: Pixel = 200;
			9871: Pixel = 205;
			9872: Pixel = 207;
			9873: Pixel = 220;
			9874: Pixel = 134;
			9875: Pixel = 73;
			9876: Pixel = 100;
			9877: Pixel = 103;
			9878: Pixel = 115;
			9879: Pixel = 120;
			9880: Pixel = 119;
			9881: Pixel = 115;
			9882: Pixel = 112;
			9883: Pixel = 114;
			9884: Pixel = 122;
			9885: Pixel = 109;
			9886: Pixel = 93;
			9887: Pixel = 97;
			9888: Pixel = 89;
			9889: Pixel = 78;
			9890: Pixel = 74;
			9891: Pixel = 81;
			9892: Pixel = 112;
			9893: Pixel = 125;
			9894: Pixel = 109;
			9895: Pixel = 81;
			9896: Pixel = 56;
			9897: Pixel = 54;
			9898: Pixel = 58;
			9899: Pixel = 74;
			9900: Pixel = 49;
			9901: Pixel = 50;
			9902: Pixel = 64;
			9903: Pixel = 176;
			9904: Pixel = 203;
			9905: Pixel = 182;
			9906: Pixel = 120;
			9907: Pixel = 148;
			9908: Pixel = 175;
			9909: Pixel = 178;
			9910: Pixel = 184;
			9911: Pixel = 157;
			9912: Pixel = 78;
			9913: Pixel = 46;
			9914: Pixel = 48;
			9915: Pixel = 54;
			9916: Pixel = 60;
			9917: Pixel = 66;
			9918: Pixel = 74;
			9919: Pixel = 58;
			9920: Pixel = 91;
			9921: Pixel = 81;
			9922: Pixel = 55;
			9923: Pixel = 89;
			9924: Pixel = 68;
			9925: Pixel = 99;
			9926: Pixel = 77;
			9927: Pixel = 92;
			9928: Pixel = 46;
			9929: Pixel = 73;
			9930: Pixel = 58;
			9931: Pixel = 66;
			9932: Pixel = 95;
			9933: Pixel = 83;
			9934: Pixel = 60;
			9935: Pixel = 84;
			9936: Pixel = 97;
			9937: Pixel = 109;
			9938: Pixel = 116;
			9939: Pixel = 121;
			9940: Pixel = 123;
			9941: Pixel = 126;
			9942: Pixel = 126;
			9943: Pixel = 127;
			9944: Pixel = 129;
			9945: Pixel = 131;
			9946: Pixel = 131;
			9947: Pixel = 134;
			9948: Pixel = 137;
			9949: Pixel = 134;
			9950: Pixel = 137;
			9951: Pixel = 139;
			9952: Pixel = 140;
			9953: Pixel = 144;
			9954: Pixel = 145;
			9955: Pixel = 143;
			9956: Pixel = 145;
			9957: Pixel = 147;
			9958: Pixel = 149;
			9959: Pixel = 148;
			9960: Pixel = 148;
			9961: Pixel = 149;
			9962: Pixel = 153;
			9963: Pixel = 155;
			9964: Pixel = 161;
			9965: Pixel = 164;
			9966: Pixel = 167;
			9967: Pixel = 174;
			9968: Pixel = 184;
			9969: Pixel = 191;
			9970: Pixel = 197;
			9971: Pixel = 202;
			9972: Pixel = 206;
			9973: Pixel = 218;
			9974: Pixel = 171;
			9975: Pixel = 84;
			9976: Pixel = 92;
			9977: Pixel = 97;
			9978: Pixel = 109;
			9979: Pixel = 122;
			9980: Pixel = 129;
			9981: Pixel = 121;
			9982: Pixel = 122;
			9983: Pixel = 134;
			9984: Pixel = 126;
			9985: Pixel = 99;
			9986: Pixel = 88;
			9987: Pixel = 79;
			9988: Pixel = 82;
			9989: Pixel = 89;
			9990: Pixel = 81;
			9991: Pixel = 100;
			9992: Pixel = 128;
			9993: Pixel = 123;
			9994: Pixel = 88;
			9995: Pixel = 57;
			9996: Pixel = 46;
			9997: Pixel = 53;
			9998: Pixel = 79;
			9999: Pixel = 100;
		endcase
	end
endmodule