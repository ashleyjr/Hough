module InHandle(
	input wire			nReset,                                                      // Common to all
	input wire			Clk,                                                        // Common to all
	output reg	[7:0]	Pixel,
	output reg			Frame,
	output reg			Line
);

	parameter COLS = 50;
	parameter ROWS = 50;
	
	reg [7:0] col;
	reg [7:0] row;
	
	always @ (posedge Clk or negedge nReset) begin
		if(!nReset) begin   
			Frame <= 0;
	    	Line  <= 0;							
			row <= ROWS-1;
			col <= COLS-1;						// Zero on first pixel	
		end else begin
			if(col == (COLS-1)) begin			// Get ready for next column
	    		Line <= 1;
				col <= 0;
				row <= row + 1;
				if(row == (ROWS-1)) begin		// Get ready for next row
					Frame <= 1;
					row <= 0;
				end
			end else begin
				Line <= 0;
				Frame <= 0;
				col = col + 1;
			end
		end
	end

	always @ (*) begin
		case(col + (row*COLS))


			0: Pixel = 159;
			1: Pixel = 157;
			2: Pixel = 153;
			3: Pixel = 158;
			4: Pixel = 173;
			5: Pixel = 150;
			6: Pixel = 97;
			7: Pixel = 101;
			8: Pixel = 106;
			9: Pixel = 105;
			10: Pixel = 112;
			11: Pixel = 123;
			12: Pixel = 128;
			13: Pixel = 130;
			14: Pixel = 129;
			15: Pixel = 131;
			16: Pixel = 133;
			17: Pixel = 132;
			18: Pixel = 132;
			19: Pixel = 133;
			20: Pixel = 132;
			21: Pixel = 130;
			22: Pixel = 130;
			23: Pixel = 131;
			24: Pixel = 132;
			25: Pixel = 131;
			26: Pixel = 129;
			27: Pixel = 129;
			28: Pixel = 128;
			29: Pixel = 126;
			30: Pixel = 114;
			31: Pixel = 113;
			32: Pixel = 151;
			33: Pixel = 156;
			34: Pixel = 152;
			35: Pixel = 154;
			36: Pixel = 152;
			37: Pixel = 155;
			38: Pixel = 151;
			39: Pixel = 178;
			40: Pixel = 223;
			41: Pixel = 136;
			42: Pixel = 108;
			43: Pixel = 123;
			44: Pixel = 121;
			45: Pixel = 123;
			46: Pixel = 122;
			47: Pixel = 124;
			48: Pixel = 127;
			49: Pixel = 116;
			50: Pixel = 156;
			51: Pixel = 156;
			52: Pixel = 154;
			53: Pixel = 162;
			54: Pixel = 169;
			55: Pixel = 145;
			56: Pixel = 95;
			57: Pixel = 99;
			58: Pixel = 106;
			59: Pixel = 102;
			60: Pixel = 111;
			61: Pixel = 122;
			62: Pixel = 126;
			63: Pixel = 129;
			64: Pixel = 130;
			65: Pixel = 130;
			66: Pixel = 132;
			67: Pixel = 132;
			68: Pixel = 131;
			69: Pixel = 131;
			70: Pixel = 132;
			71: Pixel = 131;
			72: Pixel = 129;
			73: Pixel = 132;
			74: Pixel = 132;
			75: Pixel = 130;
			76: Pixel = 129;
			77: Pixel = 127;
			78: Pixel = 128;
			79: Pixel = 127;
			80: Pixel = 118;
			81: Pixel = 106;
			82: Pixel = 135;
			83: Pixel = 159;
			84: Pixel = 159;
			85: Pixel = 160;
			86: Pixel = 156;
			87: Pixel = 154;
			88: Pixel = 151;
			89: Pixel = 152;
			90: Pixel = 210;
			91: Pixel = 193;
			92: Pixel = 107;
			93: Pixel = 118;
			94: Pixel = 121;
			95: Pixel = 122;
			96: Pixel = 124;
			97: Pixel = 135;
			98: Pixel = 94;
			99: Pixel = 44;
			100: Pixel = 156;
			101: Pixel = 157;
			102: Pixel = 160;
			103: Pixel = 165;
			104: Pixel = 162;
			105: Pixel = 146;
			106: Pixel = 95;
			107: Pixel = 99;
			108: Pixel = 106;
			109: Pixel = 103;
			110: Pixel = 111;
			111: Pixel = 121;
			112: Pixel = 126;
			113: Pixel = 128;
			114: Pixel = 129;
			115: Pixel = 130;
			116: Pixel = 130;
			117: Pixel = 130;
			118: Pixel = 131;
			119: Pixel = 131;
			120: Pixel = 126;
			121: Pixel = 128;
			122: Pixel = 128;
			123: Pixel = 130;
			124: Pixel = 132;
			125: Pixel = 130;
			126: Pixel = 127;
			127: Pixel = 126;
			128: Pixel = 126;
			129: Pixel = 127;
			130: Pixel = 122;
			131: Pixel = 107;
			132: Pixel = 124;
			133: Pixel = 158;
			134: Pixel = 162;
			135: Pixel = 160;
			136: Pixel = 157;
			137: Pixel = 154;
			138: Pixel = 154;
			139: Pixel = 145;
			140: Pixel = 168;
			141: Pixel = 227;
			142: Pixel = 151;
			143: Pixel = 107;
			144: Pixel = 124;
			145: Pixel = 121;
			146: Pixel = 136;
			147: Pixel = 92;
			148: Pixel = 40;
			149: Pixel = 50;
			150: Pixel = 159;
			151: Pixel = 161;
			152: Pixel = 167;
			153: Pixel = 163;
			154: Pixel = 161;
			155: Pixel = 145;
			156: Pixel = 92;
			157: Pixel = 99;
			158: Pixel = 104;
			159: Pixel = 102;
			160: Pixel = 110;
			161: Pixel = 120;
			162: Pixel = 124;
			163: Pixel = 126;
			164: Pixel = 126;
			165: Pixel = 128;
			166: Pixel = 128;
			167: Pixel = 129;
			168: Pixel = 129;
			169: Pixel = 127;
			170: Pixel = 121;
			171: Pixel = 120;
			172: Pixel = 118;
			173: Pixel = 119;
			174: Pixel = 127;
			175: Pixel = 131;
			176: Pixel = 127;
			177: Pixel = 126;
			178: Pixel = 125;
			179: Pixel = 126;
			180: Pixel = 120;
			181: Pixel = 110;
			182: Pixel = 123;
			183: Pixel = 150;
			184: Pixel = 158;
			185: Pixel = 157;
			186: Pixel = 156;
			187: Pixel = 155;
			188: Pixel = 156;
			189: Pixel = 152;
			190: Pixel = 142;
			191: Pixel = 200;
			192: Pixel = 216;
			193: Pixel = 116;
			194: Pixel = 113;
			195: Pixel = 133;
			196: Pixel = 89;
			197: Pixel = 41;
			198: Pixel = 53;
			199: Pixel = 50;
			200: Pixel = 160;
			201: Pixel = 166;
			202: Pixel = 156;
			203: Pixel = 156;
			204: Pixel = 163;
			205: Pixel = 145;
			206: Pixel = 91;
			207: Pixel = 98;
			208: Pixel = 105;
			209: Pixel = 102;
			210: Pixel = 111;
			211: Pixel = 120;
			212: Pixel = 123;
			213: Pixel = 125;
			214: Pixel = 127;
			215: Pixel = 128;
			216: Pixel = 126;
			217: Pixel = 129;
			218: Pixel = 128;
			219: Pixel = 132;
			220: Pixel = 135;
			221: Pixel = 146;
			222: Pixel = 153;
			223: Pixel = 145;
			224: Pixel = 132;
			225: Pixel = 119;
			226: Pixel = 125;
			227: Pixel = 130;
			228: Pixel = 126;
			229: Pixel = 126;
			230: Pixel = 120;
			231: Pixel = 110;
			232: Pixel = 120;
			233: Pixel = 144;
			234: Pixel = 151;
			235: Pixel = 155;
			236: Pixel = 153;
			237: Pixel = 154;
			238: Pixel = 151;
			239: Pixel = 146;
			240: Pixel = 139;
			241: Pixel = 158;
			242: Pixel = 229;
			243: Pixel = 170;
			244: Pixel = 109;
			245: Pixel = 90;
			246: Pixel = 39;
			247: Pixel = 55;
			248: Pixel = 53;
			249: Pixel = 45;
			250: Pixel = 165;
			251: Pixel = 161;
			252: Pixel = 130;
			253: Pixel = 156;
			254: Pixel = 167;
			255: Pixel = 147;
			256: Pixel = 89;
			257: Pixel = 94;
			258: Pixel = 102;
			259: Pixel = 103;
			260: Pixel = 112;
			261: Pixel = 121;
			262: Pixel = 124;
			263: Pixel = 125;
			264: Pixel = 127;
			265: Pixel = 128;
			266: Pixel = 133;
			267: Pixel = 129;
			268: Pixel = 134;
			269: Pixel = 145;
			270: Pixel = 153;
			271: Pixel = 169;
			272: Pixel = 178;
			273: Pixel = 182;
			274: Pixel = 187;
			275: Pixel = 169;
			276: Pixel = 127;
			277: Pixel = 119;
			278: Pixel = 127;
			279: Pixel = 123;
			280: Pixel = 116;
			281: Pixel = 107;
			282: Pixel = 120;
			283: Pixel = 144;
			284: Pixel = 145;
			285: Pixel = 151;
			286: Pixel = 150;
			287: Pixel = 147;
			288: Pixel = 145;
			289: Pixel = 141;
			290: Pixel = 141;
			291: Pixel = 136;
			292: Pixel = 186;
			293: Pixel = 238;
			294: Pixel = 114;
			295: Pixel = 33;
			296: Pixel = 53;
			297: Pixel = 52;
			298: Pixel = 48;
			299: Pixel = 48;
			300: Pixel = 173;
			301: Pixel = 132;
			302: Pixel = 104;
			303: Pixel = 162;
			304: Pixel = 167;
			305: Pixel = 146;
			306: Pixel = 84;
			307: Pixel = 89;
			308: Pixel = 99;
			309: Pixel = 100;
			310: Pixel = 108;
			311: Pixel = 115;
			312: Pixel = 119;
			313: Pixel = 123;
			314: Pixel = 125;
			315: Pixel = 126;
			316: Pixel = 124;
			317: Pixel = 123;
			318: Pixel = 130;
			319: Pixel = 133;
			320: Pixel = 142;
			321: Pixel = 156;
			322: Pixel = 171;
			323: Pixel = 181;
			324: Pixel = 187;
			325: Pixel = 199;
			326: Pixel = 192;
			327: Pixel = 141;
			328: Pixel = 103;
			329: Pixel = 115;
			330: Pixel = 114;
			331: Pixel = 103;
			332: Pixel = 118;
			333: Pixel = 149;
			334: Pixel = 146;
			335: Pixel = 144;
			336: Pixel = 148;
			337: Pixel = 142;
			338: Pixel = 144;
			339: Pixel = 142;
			340: Pixel = 142;
			341: Pixel = 139;
			342: Pixel = 157;
			343: Pixel = 195;
			344: Pixel = 60;
			345: Pixel = 44;
			346: Pixel = 54;
			347: Pixel = 48;
			348: Pixel = 50;
			349: Pixel = 43;
			350: Pixel = 161;
			351: Pixel = 95;
			352: Pixel = 102;
			353: Pixel = 163;
			354: Pixel = 168;
			355: Pixel = 143;
			356: Pixel = 83;
			357: Pixel = 91;
			358: Pixel = 100;
			359: Pixel = 100;
			360: Pixel = 107;
			361: Pixel = 114;
			362: Pixel = 118;
			363: Pixel = 121;
			364: Pixel = 128;
			365: Pixel = 114;
			366: Pixel = 112;
			367: Pixel = 123;
			368: Pixel = 127;
			369: Pixel = 133;
			370: Pixel = 135;
			371: Pixel = 148;
			372: Pixel = 170;
			373: Pixel = 185;
			374: Pixel = 188;
			375: Pixel = 189;
			376: Pixel = 196;
			377: Pixel = 208;
			378: Pixel = 175;
			379: Pixel = 101;
			380: Pixel = 106;
			381: Pixel = 101;
			382: Pixel = 117;
			383: Pixel = 153;
			384: Pixel = 153;
			385: Pixel = 124;
			386: Pixel = 128;
			387: Pixel = 148;
			388: Pixel = 144;
			389: Pixel = 143;
			390: Pixel = 143;
			391: Pixel = 148;
			392: Pixel = 149;
			393: Pixel = 59;
			394: Pixel = 39;
			395: Pixel = 52;
			396: Pixel = 48;
			397: Pixel = 52;
			398: Pixel = 52;
			399: Pixel = 82;
			400: Pixel = 122;
			401: Pixel = 81;
			402: Pixel = 108;
			403: Pixel = 161;
			404: Pixel = 168;
			405: Pixel = 142;
			406: Pixel = 85;
			407: Pixel = 91;
			408: Pixel = 100;
			409: Pixel = 101;
			410: Pixel = 107;
			411: Pixel = 115;
			412: Pixel = 120;
			413: Pixel = 123;
			414: Pixel = 115;
			415: Pixel = 111;
			416: Pixel = 119;
			417: Pixel = 118;
			418: Pixel = 125;
			419: Pixel = 135;
			420: Pixel = 138;
			421: Pixel = 145;
			422: Pixel = 169;
			423: Pixel = 180;
			424: Pixel = 183;
			425: Pixel = 200;
			426: Pixel = 206;
			427: Pixel = 206;
			428: Pixel = 228;
			429: Pixel = 167;
			430: Pixel = 79;
			431: Pixel = 96;
			432: Pixel = 115;
			433: Pixel = 152;
			434: Pixel = 157;
			435: Pixel = 115;
			436: Pixel = 77;
			437: Pixel = 143;
			438: Pixel = 146;
			439: Pixel = 143;
			440: Pixel = 142;
			441: Pixel = 155;
			442: Pixel = 87;
			443: Pixel = 37;
			444: Pixel = 55;
			445: Pixel = 49;
			446: Pixel = 49;
			447: Pixel = 55;
			448: Pixel = 92;
			449: Pixel = 147;
			450: Pixel = 91;
			451: Pixel = 87;
			452: Pixel = 106;
			453: Pixel = 158;
			454: Pixel = 168;
			455: Pixel = 142;
			456: Pixel = 85;
			457: Pixel = 92;
			458: Pixel = 100;
			459: Pixel = 100;
			460: Pixel = 106;
			461: Pixel = 116;
			462: Pixel = 120;
			463: Pixel = 120;
			464: Pixel = 110;
			465: Pixel = 115;
			466: Pixel = 115;
			467: Pixel = 121;
			468: Pixel = 133;
			469: Pixel = 139;
			470: Pixel = 142;
			471: Pixel = 140;
			472: Pixel = 157;
			473: Pixel = 180;
			474: Pixel = 201;
			475: Pixel = 203;
			476: Pixel = 200;
			477: Pixel = 203;
			478: Pixel = 206;
			479: Pixel = 222;
			480: Pixel = 150;
			481: Pixel = 74;
			482: Pixel = 114;
			483: Pixel = 153;
			484: Pixel = 157;
			485: Pixel = 122;
			486: Pixel = 46;
			487: Pixel = 112;
			488: Pixel = 150;
			489: Pixel = 137;
			490: Pixel = 154;
			491: Pixel = 119;
			492: Pixel = 38;
			493: Pixel = 55;
			494: Pixel = 49;
			495: Pixel = 51;
			496: Pixel = 48;
			497: Pixel = 82;
			498: Pixel = 145;
			499: Pixel = 155;
			500: Pixel = 91;
			501: Pixel = 88;
			502: Pixel = 107;
			503: Pixel = 157;
			504: Pixel = 166;
			505: Pixel = 144;
			506: Pixel = 86;
			507: Pixel = 89;
			508: Pixel = 100;
			509: Pixel = 100;
			510: Pixel = 107;
			511: Pixel = 113;
			512: Pixel = 128;
			513: Pixel = 114;
			514: Pixel = 108;
			515: Pixel = 113;
			516: Pixel = 119;
			517: Pixel = 133;
			518: Pixel = 138;
			519: Pixel = 140;
			520: Pixel = 125;
			521: Pixel = 142;
			522: Pixel = 181;
			523: Pixel = 194;
			524: Pixel = 190;
			525: Pixel = 195;
			526: Pixel = 203;
			527: Pixel = 204;
			528: Pixel = 204;
			529: Pixel = 204;
			530: Pixel = 231;
			531: Pixel = 131;
			532: Pixel = 95;
			533: Pixel = 154;
			534: Pixel = 156;
			535: Pixel = 125;
			536: Pixel = 48;
			537: Pixel = 49;
			538: Pixel = 131;
			539: Pixel = 154;
			540: Pixel = 139;
			541: Pixel = 55;
			542: Pixel = 46;
			543: Pixel = 55;
			544: Pixel = 51;
			545: Pixel = 47;
			546: Pixel = 61;
			547: Pixel = 135;
			548: Pixel = 151;
			549: Pixel = 163;
			550: Pixel = 91;
			551: Pixel = 86;
			552: Pixel = 103;
			553: Pixel = 157;
			554: Pixel = 166;
			555: Pixel = 144;
			556: Pixel = 82;
			557: Pixel = 86;
			558: Pixel = 98;
			559: Pixel = 99;
			560: Pixel = 107;
			561: Pixel = 108;
			562: Pixel = 148;
			563: Pixel = 109;
			564: Pixel = 109;
			565: Pixel = 115;
			566: Pixel = 125;
			567: Pixel = 131;
			568: Pixel = 133;
			569: Pixel = 121;
			570: Pixel = 144;
			571: Pixel = 179;
			572: Pixel = 182;
			573: Pixel = 181;
			574: Pixel = 192;
			575: Pixel = 196;
			576: Pixel = 197;
			577: Pixel = 200;
			578: Pixel = 202;
			579: Pixel = 204;
			580: Pixel = 212;
			581: Pixel = 205;
			582: Pixel = 101;
			583: Pixel = 148;
			584: Pixel = 159;
			585: Pixel = 125;
			586: Pixel = 35;
			587: Pixel = 77;
			588: Pixel = 186;
			589: Pixel = 226;
			590: Pixel = 158;
			591: Pixel = 35;
			592: Pixel = 57;
			593: Pixel = 52;
			594: Pixel = 53;
			595: Pixel = 48;
			596: Pixel = 119;
			597: Pixel = 153;
			598: Pixel = 159;
			599: Pixel = 158;
			600: Pixel = 94;
			601: Pixel = 94;
			602: Pixel = 105;
			603: Pixel = 157;
			604: Pixel = 169;
			605: Pixel = 145;
			606: Pixel = 82;
			607: Pixel = 88;
			608: Pixel = 101;
			609: Pixel = 100;
			610: Pixel = 106;
			611: Pixel = 118;
			612: Pixel = 160;
			613: Pixel = 100;
			614: Pixel = 108;
			615: Pixel = 119;
			616: Pixel = 124;
			617: Pixel = 126;
			618: Pixel = 120;
			619: Pixel = 147;
			620: Pixel = 172;
			621: Pixel = 171;
			622: Pixel = 178;
			623: Pixel = 185;
			624: Pixel = 184;
			625: Pixel = 186;
			626: Pixel = 195;
			627: Pixel = 198;
			628: Pixel = 198;
			629: Pixel = 198;
			630: Pixel = 202;
			631: Pixel = 213;
			632: Pixel = 169;
			633: Pixel = 142;
			634: Pixel = 157;
			635: Pixel = 108;
			636: Pixel = 111;
			637: Pixel = 201;
			638: Pixel = 210;
			639: Pixel = 216;
			640: Pixel = 195;
			641: Pixel = 47;
			642: Pixel = 51;
			643: Pixel = 49;
			644: Pixel = 41;
			645: Pixel = 90;
			646: Pixel = 155;
			647: Pixel = 156;
			648: Pixel = 158;
			649: Pixel = 156;
			650: Pixel = 100;
			651: Pixel = 97;
			652: Pixel = 110;
			653: Pixel = 157;
			654: Pixel = 172;
			655: Pixel = 150;
			656: Pixel = 85;
			657: Pixel = 91;
			658: Pixel = 102;
			659: Pixel = 101;
			660: Pixel = 102;
			661: Pixel = 125;
			662: Pixel = 158;
			663: Pixel = 98;
			664: Pixel = 105;
			665: Pixel = 114;
			666: Pixel = 121;
			667: Pixel = 121;
			668: Pixel = 143;
			669: Pixel = 152;
			670: Pixel = 158;
			671: Pixel = 174;
			672: Pixel = 176;
			673: Pixel = 175;
			674: Pixel = 175;
			675: Pixel = 182;
			676: Pixel = 187;
			677: Pixel = 192;
			678: Pixel = 184;
			679: Pixel = 189;
			680: Pixel = 199;
			681: Pixel = 195;
			682: Pixel = 205;
			683: Pixel = 168;
			684: Pixel = 155;
			685: Pixel = 181;
			686: Pixel = 209;
			687: Pixel = 205;
			688: Pixel = 200;
			689: Pixel = 218;
			690: Pixel = 179;
			691: Pixel = 43;
			692: Pixel = 51;
			693: Pixel = 47;
			694: Pixel = 58;
			695: Pixel = 139;
			696: Pixel = 158;
			697: Pixel = 158;
			698: Pixel = 155;
			699: Pixel = 154;
			700: Pixel = 99;
			701: Pixel = 96;
			702: Pixel = 111;
			703: Pixel = 159;
			704: Pixel = 176;
			705: Pixel = 152;
			706: Pixel = 85;
			707: Pixel = 90;
			708: Pixel = 100;
			709: Pixel = 99;
			710: Pixel = 96;
			711: Pixel = 133;
			712: Pixel = 170;
			713: Pixel = 110;
			714: Pixel = 106;
			715: Pixel = 114;
			716: Pixel = 119;
			717: Pixel = 140;
			718: Pixel = 143;
			719: Pixel = 143;
			720: Pixel = 155;
			721: Pixel = 166;
			722: Pixel = 167;
			723: Pixel = 170;
			724: Pixel = 175;
			725: Pixel = 173;
			726: Pixel = 179;
			727: Pixel = 179;
			728: Pixel = 184;
			729: Pixel = 189;
			730: Pixel = 183;
			731: Pixel = 180;
			732: Pixel = 177;
			733: Pixel = 188;
			734: Pixel = 198;
			735: Pixel = 205;
			736: Pixel = 199;
			737: Pixel = 201;
			738: Pixel = 192;
			739: Pixel = 220;
			740: Pixel = 144;
			741: Pixel = 35;
			742: Pixel = 52;
			743: Pixel = 45;
			744: Pixel = 114;
			745: Pixel = 156;
			746: Pixel = 159;
			747: Pixel = 158;
			748: Pixel = 156;
			749: Pixel = 155;
			750: Pixel = 97;
			751: Pixel = 93;
			752: Pixel = 109;
			753: Pixel = 161;
			754: Pixel = 175;
			755: Pixel = 152;
			756: Pixel = 87;
			757: Pixel = 92;
			758: Pixel = 100;
			759: Pixel = 100;
			760: Pixel = 94;
			761: Pixel = 135;
			762: Pixel = 177;
			763: Pixel = 132;
			764: Pixel = 103;
			765: Pixel = 112;
			766: Pixel = 134;
			767: Pixel = 134;
			768: Pixel = 138;
			769: Pixel = 147;
			770: Pixel = 147;
			771: Pixel = 158;
			772: Pixel = 169;
			773: Pixel = 168;
			774: Pixel = 168;
			775: Pixel = 163;
			776: Pixel = 166;
			777: Pixel = 175;
			778: Pixel = 180;
			779: Pixel = 173;
			780: Pixel = 169;
			781: Pixel = 173;
			782: Pixel = 190;
			783: Pixel = 197;
			784: Pixel = 196;
			785: Pixel = 196;
			786: Pixel = 199;
			787: Pixel = 203;
			788: Pixel = 165;
			789: Pixel = 183;
			790: Pixel = 87;
			791: Pixel = 41;
			792: Pixel = 45;
			793: Pixel = 77;
			794: Pixel = 148;
			795: Pixel = 157;
			796: Pixel = 160;
			797: Pixel = 158;
			798: Pixel = 157;
			799: Pixel = 157;
			800: Pixel = 96;
			801: Pixel = 94;
			802: Pixel = 113;
			803: Pixel = 161;
			804: Pixel = 174;
			805: Pixel = 154;
			806: Pixel = 86;
			807: Pixel = 90;
			808: Pixel = 98;
			809: Pixel = 99;
			810: Pixel = 89;
			811: Pixel = 139;
			812: Pixel = 186;
			813: Pixel = 147;
			814: Pixel = 116;
			815: Pixel = 126;
			816: Pixel = 130;
			817: Pixel = 133;
			818: Pixel = 138;
			819: Pixel = 137;
			820: Pixel = 148;
			821: Pixel = 145;
			822: Pixel = 141;
			823: Pixel = 145;
			824: Pixel = 148;
			825: Pixel = 160;
			826: Pixel = 165;
			827: Pixel = 161;
			828: Pixel = 152;
			829: Pixel = 161;
			830: Pixel = 178;
			831: Pixel = 193;
			832: Pixel = 193;
			833: Pixel = 193;
			834: Pixel = 196;
			835: Pixel = 204;
			836: Pixel = 218;
			837: Pixel = 175;
			838: Pixel = 131;
			839: Pixel = 162;
			840: Pixel = 48;
			841: Pixel = 50;
			842: Pixel = 51;
			843: Pixel = 124;
			844: Pixel = 157;
			845: Pixel = 158;
			846: Pixel = 156;
			847: Pixel = 156;
			848: Pixel = 156;
			849: Pixel = 155;
			850: Pixel = 99;
			851: Pixel = 98;
			852: Pixel = 118;
			853: Pixel = 162;
			854: Pixel = 176;
			855: Pixel = 156;
			856: Pixel = 84;
			857: Pixel = 89;
			858: Pixel = 99;
			859: Pixel = 101;
			860: Pixel = 88;
			861: Pixel = 136;
			862: Pixel = 201;
			863: Pixel = 146;
			864: Pixel = 125;
			865: Pixel = 116;
			866: Pixel = 129;
			867: Pixel = 134;
			868: Pixel = 128;
			869: Pixel = 136;
			870: Pixel = 138;
			871: Pixel = 126;
			872: Pixel = 94;
			873: Pixel = 115;
			874: Pixel = 120;
			875: Pixel = 100;
			876: Pixel = 90;
			877: Pixel = 59;
			878: Pixel = 123;
			879: Pixel = 186;
			880: Pixel = 195;
			881: Pixel = 195;
			882: Pixel = 191;
			883: Pixel = 200;
			884: Pixel = 210;
			885: Pixel = 192;
			886: Pixel = 148;
			887: Pixel = 96;
			888: Pixel = 154;
			889: Pixel = 108;
			890: Pixel = 37;
			891: Pixel = 46;
			892: Pixel = 74;
			893: Pixel = 150;
			894: Pixel = 158;
			895: Pixel = 159;
			896: Pixel = 156;
			897: Pixel = 154;
			898: Pixel = 154;
			899: Pixel = 153;
			900: Pixel = 103;
			901: Pixel = 98;
			902: Pixel = 118;
			903: Pixel = 162;
			904: Pixel = 175;
			905: Pixel = 156;
			906: Pixel = 86;
			907: Pixel = 88;
			908: Pixel = 99;
			909: Pixel = 100;
			910: Pixel = 93;
			911: Pixel = 113;
			912: Pixel = 203;
			913: Pixel = 146;
			914: Pixel = 123;
			915: Pixel = 120;
			916: Pixel = 131;
			917: Pixel = 125;
			918: Pixel = 132;
			919: Pixel = 134;
			920: Pixel = 114;
			921: Pixel = 92;
			922: Pixel = 66;
			923: Pixel = 85;
			924: Pixel = 87;
			925: Pixel = 75;
			926: Pixel = 50;
			927: Pixel = 104;
			928: Pixel = 177;
			929: Pixel = 190;
			930: Pixel = 190;
			931: Pixel = 189;
			932: Pixel = 198;
			933: Pixel = 192;
			934: Pixel = 157;
			935: Pixel = 115;
			936: Pixel = 109;
			937: Pixel = 170;
			938: Pixel = 111;
			939: Pixel = 40;
			940: Pixel = 51;
			941: Pixel = 48;
			942: Pixel = 113;
			943: Pixel = 160;
			944: Pixel = 162;
			945: Pixel = 160;
			946: Pixel = 158;
			947: Pixel = 155;
			948: Pixel = 154;
			949: Pixel = 153;
			950: Pixel = 106;
			951: Pixel = 99;
			952: Pixel = 114;
			953: Pixel = 161;
			954: Pixel = 174;
			955: Pixel = 156;
			956: Pixel = 86;
			957: Pixel = 87;
			958: Pixel = 98;
			959: Pixel = 97;
			960: Pixel = 100;
			961: Pixel = 95;
			962: Pixel = 182;
			963: Pixel = 177;
			964: Pixel = 125;
			965: Pixel = 127;
			966: Pixel = 121;
			967: Pixel = 126;
			968: Pixel = 124;
			969: Pixel = 99;
			970: Pixel = 73;
			971: Pixel = 57;
			972: Pixel = 58;
			973: Pixel = 71;
			974: Pixel = 80;
			975: Pixel = 72;
			976: Pixel = 122;
			977: Pixel = 189;
			978: Pixel = 186;
			979: Pixel = 178;
			980: Pixel = 178;
			981: Pixel = 192;
			982: Pixel = 171;
			983: Pixel = 96;
			984: Pixel = 107;
			985: Pixel = 155;
			986: Pixel = 189;
			987: Pixel = 107;
			988: Pixel = 36;
			989: Pixel = 56;
			990: Pixel = 46;
			991: Pixel = 64;
			992: Pixel = 141;
			993: Pixel = 163;
			994: Pixel = 164;
			995: Pixel = 162;
			996: Pixel = 159;
			997: Pixel = 157;
			998: Pixel = 155;
			999: Pixel = 152;
			1000: Pixel = 107;
			1001: Pixel = 98;
			1002: Pixel = 106;
			1003: Pixel = 160;
			1004: Pixel = 176;
			1005: Pixel = 158;
			1006: Pixel = 85;
			1007: Pixel = 85;
			1008: Pixel = 98;
			1009: Pixel = 96;
			1010: Pixel = 104;
			1011: Pixel = 99;
			1012: Pixel = 135;
			1013: Pixel = 198;
			1014: Pixel = 126;
			1015: Pixel = 118;
			1016: Pixel = 127;
			1017: Pixel = 126;
			1018: Pixel = 91;
			1019: Pixel = 74;
			1020: Pixel = 62;
			1021: Pixel = 69;
			1022: Pixel = 60;
			1023: Pixel = 53;
			1024: Pixel = 63;
			1025: Pixel = 108;
			1026: Pixel = 170;
			1027: Pixel = 186;
			1028: Pixel = 175;
			1029: Pixel = 174;
			1030: Pixel = 181;
			1031: Pixel = 194;
			1032: Pixel = 177;
			1033: Pixel = 89;
			1034: Pixel = 102;
			1035: Pixel = 151;
			1036: Pixel = 86;
			1037: Pixel = 33;
			1038: Pixel = 58;
			1039: Pixel = 51;
			1040: Pixel = 45;
			1041: Pixel = 93;
			1042: Pixel = 146;
			1043: Pixel = 168;
			1044: Pixel = 163;
			1045: Pixel = 162;
			1046: Pixel = 160;
			1047: Pixel = 159;
			1048: Pixel = 156;
			1049: Pixel = 153;
			1050: Pixel = 105;
			1051: Pixel = 98;
			1052: Pixel = 103;
			1053: Pixel = 158;
			1054: Pixel = 176;
			1055: Pixel = 159;
			1056: Pixel = 86;
			1057: Pixel = 86;
			1058: Pixel = 101;
			1059: Pixel = 98;
			1060: Pixel = 105;
			1061: Pixel = 108;
			1062: Pixel = 128;
			1063: Pixel = 184;
			1064: Pixel = 108;
			1065: Pixel = 120;
			1066: Pixel = 124;
			1067: Pixel = 87;
			1068: Pixel = 54;
			1069: Pixel = 54;
			1070: Pixel = 68;
			1071: Pixel = 74;
			1072: Pixel = 67;
			1073: Pixel = 41;
			1074: Pixel = 111;
			1075: Pixel = 150;
			1076: Pixel = 184;
			1077: Pixel = 169;
			1078: Pixel = 167;
			1079: Pixel = 173;
			1080: Pixel = 195;
			1081: Pixel = 200;
			1082: Pixel = 208;
			1083: Pixel = 108;
			1084: Pixel = 57;
			1085: Pixel = 134;
			1086: Pixel = 50;
			1087: Pixel = 51;
			1088: Pixel = 61;
			1089: Pixel = 47;
			1090: Pixel = 54;
			1091: Pixel = 125;
			1092: Pixel = 150;
			1093: Pixel = 160;
			1094: Pixel = 162;
			1095: Pixel = 162;
			1096: Pixel = 162;
			1097: Pixel = 159;
			1098: Pixel = 157;
			1099: Pixel = 153;
			1100: Pixel = 104;
			1101: Pixel = 97;
			1102: Pixel = 103;
			1103: Pixel = 158;
			1104: Pixel = 177;
			1105: Pixel = 159;
			1106: Pixel = 90;
			1107: Pixel = 89;
			1108: Pixel = 103;
			1109: Pixel = 100;
			1110: Pixel = 109;
			1111: Pixel = 117;
			1112: Pixel = 119;
			1113: Pixel = 150;
			1114: Pixel = 115;
			1115: Pixel = 127;
			1116: Pixel = 77;
			1117: Pixel = 52;
			1118: Pixel = 60;
			1119: Pixel = 52;
			1120: Pixel = 56;
			1121: Pixel = 77;
			1122: Pixel = 65;
			1123: Pixel = 108;
			1124: Pixel = 179;
			1125: Pixel = 165;
			1126: Pixel = 181;
			1127: Pixel = 164;
			1128: Pixel = 161;
			1129: Pixel = 185;
			1130: Pixel = 199;
			1131: Pixel = 203;
			1132: Pixel = 216;
			1133: Pixel = 146;
			1134: Pixel = 41;
			1135: Pixel = 119;
			1136: Pixel = 66;
			1137: Pixel = 54;
			1138: Pixel = 59;
			1139: Pixel = 43;
			1140: Pixel = 79;
			1141: Pixel = 149;
			1142: Pixel = 159;
			1143: Pixel = 152;
			1144: Pixel = 151;
			1145: Pixel = 151;
			1146: Pixel = 155;
			1147: Pixel = 156;
			1148: Pixel = 155;
			1149: Pixel = 153;
			1150: Pixel = 102;
			1151: Pixel = 95;
			1152: Pixel = 102;
			1153: Pixel = 159;
			1154: Pixel = 178;
			1155: Pixel = 159;
			1156: Pixel = 89;
			1157: Pixel = 90;
			1158: Pixel = 103;
			1159: Pixel = 102;
			1160: Pixel = 109;
			1161: Pixel = 117;
			1162: Pixel = 119;
			1163: Pixel = 112;
			1164: Pixel = 136;
			1165: Pixel = 93;
			1166: Pixel = 59;
			1167: Pixel = 57;
			1168: Pixel = 63;
			1169: Pixel = 51;
			1170: Pixel = 64;
			1171: Pixel = 53;
			1172: Pixel = 92;
			1173: Pixel = 163;
			1174: Pixel = 178;
			1175: Pixel = 177;
			1176: Pixel = 148;
			1177: Pixel = 157;
			1178: Pixel = 177;
			1179: Pixel = 183;
			1180: Pixel = 195;
			1181: Pixel = 198;
			1182: Pixel = 221;
			1183: Pixel = 172;
			1184: Pixel = 42;
			1185: Pixel = 102;
			1186: Pixel = 80;
			1187: Pixel = 56;
			1188: Pixel = 56;
			1189: Pixel = 47;
			1190: Pixel = 111;
			1191: Pixel = 156;
			1192: Pixel = 162;
			1193: Pixel = 161;
			1194: Pixel = 161;
			1195: Pixel = 151;
			1196: Pixel = 146;
			1197: Pixel = 143;
			1198: Pixel = 145;
			1199: Pixel = 148;
			1200: Pixel = 102;
			1201: Pixel = 99;
			1202: Pixel = 101;
			1203: Pixel = 158;
			1204: Pixel = 179;
			1205: Pixel = 162;
			1206: Pixel = 90;
			1207: Pixel = 89;
			1208: Pixel = 103;
			1209: Pixel = 100;
			1210: Pixel = 103;
			1211: Pixel = 126;
			1212: Pixel = 136;
			1213: Pixel = 89;
			1214: Pixel = 105;
			1215: Pixel = 70;
			1216: Pixel = 74;
			1217: Pixel = 59;
			1218: Pixel = 58;
			1219: Pixel = 50;
			1220: Pixel = 59;
			1221: Pixel = 71;
			1222: Pixel = 157;
			1223: Pixel = 185;
			1224: Pixel = 172;
			1225: Pixel = 136;
			1226: Pixel = 111;
			1227: Pixel = 98;
			1228: Pixel = 137;
			1229: Pixel = 172;
			1230: Pixel = 187;
			1231: Pixel = 197;
			1232: Pixel = 152;
			1233: Pixel = 108;
			1234: Pixel = 50;
			1235: Pixel = 91;
			1236: Pixel = 94;
			1237: Pixel = 56;
			1238: Pixel = 50;
			1239: Pixel = 61;
			1240: Pixel = 132;
			1241: Pixel = 158;
			1242: Pixel = 157;
			1243: Pixel = 156;
			1244: Pixel = 159;
			1245: Pixel = 155;
			1246: Pixel = 154;
			1247: Pixel = 153;
			1248: Pixel = 145;
			1249: Pixel = 137;
			1250: Pixel = 99;
			1251: Pixel = 92;
			1252: Pixel = 93;
			1253: Pixel = 158;
			1254: Pixel = 179;
			1255: Pixel = 161;
			1256: Pixel = 89;
			1257: Pixel = 87;
			1258: Pixel = 102;
			1259: Pixel = 93;
			1260: Pixel = 121;
			1261: Pixel = 158;
			1262: Pixel = 141;
			1263: Pixel = 78;
			1264: Pixel = 65;
			1265: Pixel = 86;
			1266: Pixel = 69;
			1267: Pixel = 58;
			1268: Pixel = 57;
			1269: Pixel = 63;
			1270: Pixel = 40;
			1271: Pixel = 128;
			1272: Pixel = 195;
			1273: Pixel = 176;
			1274: Pixel = 75;
			1275: Pixel = 49;
			1276: Pixel = 86;
			1277: Pixel = 84;
			1278: Pixel = 113;
			1279: Pixel = 149;
			1280: Pixel = 199;
			1281: Pixel = 124;
			1282: Pixel = 66;
			1283: Pixel = 67;
			1284: Pixel = 44;
			1285: Pixel = 87;
			1286: Pixel = 103;
			1287: Pixel = 53;
			1288: Pixel = 44;
			1289: Pixel = 81;
			1290: Pixel = 149;
			1291: Pixel = 157;
			1292: Pixel = 153;
			1293: Pixel = 153;
			1294: Pixel = 154;
			1295: Pixel = 153;
			1296: Pixel = 152;
			1297: Pixel = 152;
			1298: Pixel = 142;
			1299: Pixel = 133;
			1300: Pixel = 100;
			1301: Pixel = 89;
			1302: Pixel = 87;
			1303: Pixel = 158;
			1304: Pixel = 183;
			1305: Pixel = 163;
			1306: Pixel = 92;
			1307: Pixel = 95;
			1308: Pixel = 106;
			1309: Pixel = 78;
			1310: Pixel = 133;
			1311: Pixel = 162;
			1312: Pixel = 70;
			1313: Pixel = 62;
			1314: Pixel = 65;
			1315: Pixel = 94;
			1316: Pixel = 77;
			1317: Pixel = 46;
			1318: Pixel = 55;
			1319: Pixel = 37;
			1320: Pixel = 81;
			1321: Pixel = 175;
			1322: Pixel = 185;
			1323: Pixel = 126;
			1324: Pixel = 92;
			1325: Pixel = 87;
			1326: Pixel = 159;
			1327: Pixel = 156;
			1328: Pixel = 108;
			1329: Pixel = 148;
			1330: Pixel = 194;
			1331: Pixel = 96;
			1332: Pixel = 126;
			1333: Pixel = 83;
			1334: Pixel = 36;
			1335: Pixel = 88;
			1336: Pixel = 112;
			1337: Pixel = 52;
			1338: Pixel = 46;
			1339: Pixel = 109;
			1340: Pixel = 157;
			1341: Pixel = 154;
			1342: Pixel = 151;
			1343: Pixel = 153;
			1344: Pixel = 152;
			1345: Pixel = 150;
			1346: Pixel = 145;
			1347: Pixel = 135;
			1348: Pixel = 137;
			1349: Pixel = 157;
			1350: Pixel = 101;
			1351: Pixel = 85;
			1352: Pixel = 82;
			1353: Pixel = 157;
			1354: Pixel = 184;
			1355: Pixel = 167;
			1356: Pixel = 96;
			1357: Pixel = 98;
			1358: Pixel = 111;
			1359: Pixel = 125;
			1360: Pixel = 114;
			1361: Pixel = 58;
			1362: Pixel = 86;
			1363: Pixel = 83;
			1364: Pixel = 63;
			1365: Pixel = 108;
			1366: Pixel = 97;
			1367: Pixel = 42;
			1368: Pixel = 46;
			1369: Pixel = 47;
			1370: Pixel = 145;
			1371: Pixel = 185;
			1372: Pixel = 116;
			1373: Pixel = 139;
			1374: Pixel = 156;
			1375: Pixel = 143;
			1376: Pixel = 149;
			1377: Pixel = 159;
			1378: Pixel = 130;
			1379: Pixel = 139;
			1380: Pixel = 201;
			1381: Pixel = 159;
			1382: Pixel = 124;
			1383: Pixel = 89;
			1384: Pixel = 49;
			1385: Pixel = 84;
			1386: Pixel = 119;
			1387: Pixel = 44;
			1388: Pixel = 57;
			1389: Pixel = 131;
			1390: Pixel = 156;
			1391: Pixel = 152;
			1392: Pixel = 151;
			1393: Pixel = 151;
			1394: Pixel = 149;
			1395: Pixel = 143;
			1396: Pixel = 134;
			1397: Pixel = 160;
			1398: Pixel = 186;
			1399: Pixel = 191;
			1400: Pixel = 89;
			1401: Pixel = 75;
			1402: Pixel = 74;
			1403: Pixel = 155;
			1404: Pixel = 183;
			1405: Pixel = 167;
			1406: Pixel = 94;
			1407: Pixel = 95;
			1408: Pixel = 126;
			1409: Pixel = 121;
			1410: Pixel = 71;
			1411: Pixel = 72;
			1412: Pixel = 106;
			1413: Pixel = 56;
			1414: Pixel = 59;
			1415: Pixel = 90;
			1416: Pixel = 92;
			1417: Pixel = 60;
			1418: Pixel = 37;
			1419: Pixel = 97;
			1420: Pixel = 186;
			1421: Pixel = 103;
			1422: Pixel = 110;
			1423: Pixel = 146;
			1424: Pixel = 165;
			1425: Pixel = 175;
			1426: Pixel = 175;
			1427: Pixel = 163;
			1428: Pixel = 139;
			1429: Pixel = 133;
			1430: Pixel = 201;
			1431: Pixel = 173;
			1432: Pixel = 138;
			1433: Pixel = 116;
			1434: Pixel = 53;
			1435: Pixel = 78;
			1436: Pixel = 120;
			1437: Pixel = 37;
			1438: Pixel = 73;
			1439: Pixel = 147;
			1440: Pixel = 156;
			1441: Pixel = 151;
			1442: Pixel = 150;
			1443: Pixel = 148;
			1444: Pixel = 145;
			1445: Pixel = 133;
			1446: Pixel = 164;
			1447: Pixel = 200;
			1448: Pixel = 192;
			1449: Pixel = 192;
			1450: Pixel = 78;
			1451: Pixel = 68;
			1452: Pixel = 72;
			1453: Pixel = 154;
			1454: Pixel = 179;
			1455: Pixel = 164;
			1456: Pixel = 93;
			1457: Pixel = 100;
			1458: Pixel = 118;
			1459: Pixel = 95;
			1460: Pixel = 82;
			1461: Pixel = 83;
			1462: Pixel = 96;
			1463: Pixel = 49;
			1464: Pixel = 49;
			1465: Pixel = 49;
			1466: Pixel = 97;
			1467: Pixel = 97;
			1468: Pixel = 38;
			1469: Pixel = 165;
			1470: Pixel = 129;
			1471: Pixel = 56;
			1472: Pixel = 127;
			1473: Pixel = 138;
			1474: Pixel = 157;
			1475: Pixel = 174;
			1476: Pixel = 174;
			1477: Pixel = 156;
			1478: Pixel = 136;
			1479: Pixel = 127;
			1480: Pixel = 194;
			1481: Pixel = 173;
			1482: Pixel = 142;
			1483: Pixel = 109;
			1484: Pixel = 51;
			1485: Pixel = 71;
			1486: Pixel = 125;
			1487: Pixel = 42;
			1488: Pixel = 98;
			1489: Pixel = 159;
			1490: Pixel = 155;
			1491: Pixel = 150;
			1492: Pixel = 147;
			1493: Pixel = 145;
			1494: Pixel = 137;
			1495: Pixel = 147;
			1496: Pixel = 195;
			1497: Pixel = 192;
			1498: Pixel = 200;
			1499: Pixel = 203;
			1500: Pixel = 80;
			1501: Pixel = 65;
			1502: Pixel = 62;
			1503: Pixel = 153;
			1504: Pixel = 178;
			1505: Pixel = 164;
			1506: Pixel = 91;
			1507: Pixel = 111;
			1508: Pixel = 112;
			1509: Pixel = 90;
			1510: Pixel = 83;
			1511: Pixel = 91;
			1512: Pixel = 104;
			1513: Pixel = 51;
			1514: Pixel = 46;
			1515: Pixel = 86;
			1516: Pixel = 112;
			1517: Pixel = 61;
			1518: Pixel = 93;
			1519: Pixel = 161;
			1520: Pixel = 45;
			1521: Pixel = 74;
			1522: Pixel = 119;
			1523: Pixel = 136;
			1524: Pixel = 149;
			1525: Pixel = 158;
			1526: Pixel = 165;
			1527: Pixel = 145;
			1528: Pixel = 128;
			1529: Pixel = 125;
			1530: Pixel = 187;
			1531: Pixel = 177;
			1532: Pixel = 140;
			1533: Pixel = 89;
			1534: Pixel = 51;
			1535: Pixel = 63;
			1536: Pixel = 128;
			1537: Pixel = 53;
			1538: Pixel = 122;
			1539: Pixel = 160;
			1540: Pixel = 152;
			1541: Pixel = 150;
			1542: Pixel = 148;
			1543: Pixel = 144;
			1544: Pixel = 134;
			1545: Pixel = 180;
			1546: Pixel = 196;
			1547: Pixel = 200;
			1548: Pixel = 207;
			1549: Pixel = 205;
			1550: Pixel = 82;
			1551: Pixel = 67;
			1552: Pixel = 71;
			1553: Pixel = 155;
			1554: Pixel = 178;
			1555: Pixel = 166;
			1556: Pixel = 98;
			1557: Pixel = 100;
			1558: Pixel = 97;
			1559: Pixel = 84;
			1560: Pixel = 82;
			1561: Pixel = 84;
			1562: Pixel = 112;
			1563: Pixel = 64;
			1564: Pixel = 52;
			1565: Pixel = 75;
			1566: Pixel = 56;
			1567: Pixel = 63;
			1568: Pixel = 178;
			1569: Pixel = 77;
			1570: Pixel = 40;
			1571: Pixel = 89;
			1572: Pixel = 117;
			1573: Pixel = 133;
			1574: Pixel = 145;
			1575: Pixel = 152;
			1576: Pixel = 158;
			1577: Pixel = 143;
			1578: Pixel = 120;
			1579: Pixel = 108;
			1580: Pixel = 162;
			1581: Pixel = 166;
			1582: Pixel = 131;
			1583: Pixel = 59;
			1584: Pixel = 57;
			1585: Pixel = 54;
			1586: Pixel = 122;
			1587: Pixel = 80;
			1588: Pixel = 142;
			1589: Pixel = 156;
			1590: Pixel = 150;
			1591: Pixel = 149;
			1592: Pixel = 148;
			1593: Pixel = 140;
			1594: Pixel = 147;
			1595: Pixel = 195;
			1596: Pixel = 199;
			1597: Pixel = 207;
			1598: Pixel = 207;
			1599: Pixel = 207;
			1600: Pixel = 79;
			1601: Pixel = 68;
			1602: Pixel = 95;
			1603: Pixel = 160;
			1604: Pixel = 174;
			1605: Pixel = 169;
			1606: Pixel = 93;
			1607: Pixel = 97;
			1608: Pixel = 100;
			1609: Pixel = 76;
			1610: Pixel = 73;
			1611: Pixel = 77;
			1612: Pixel = 114;
			1613: Pixel = 96;
			1614: Pixel = 77;
			1615: Pixel = 54;
			1616: Pixel = 119;
			1617: Pixel = 134;
			1618: Pixel = 107;
			1619: Pixel = 43;
			1620: Pixel = 57;
			1621: Pixel = 96;
			1622: Pixel = 120;
			1623: Pixel = 131;
			1624: Pixel = 141;
			1625: Pixel = 148;
			1626: Pixel = 157;
			1627: Pixel = 155;
			1628: Pixel = 142;
			1629: Pixel = 160;
			1630: Pixel = 184;
			1631: Pixel = 157;
			1632: Pixel = 105;
			1633: Pixel = 43;
			1634: Pixel = 72;
			1635: Pixel = 55;
			1636: Pixel = 105;
			1637: Pixel = 116;
			1638: Pixel = 150;
			1639: Pixel = 154;
			1640: Pixel = 149;
			1641: Pixel = 147;
			1642: Pixel = 146;
			1643: Pixel = 136;
			1644: Pixel = 160;
			1645: Pixel = 200;
			1646: Pixel = 206;
			1647: Pixel = 207;
			1648: Pixel = 209;
			1649: Pixel = 209;
			1650: Pixel = 69;
			1651: Pixel = 63;
			1652: Pixel = 94;
			1653: Pixel = 161;
			1654: Pixel = 176;
			1655: Pixel = 170;
			1656: Pixel = 92;
			1657: Pixel = 105;
			1658: Pixel = 98;
			1659: Pixel = 78;
			1660: Pixel = 61;
			1661: Pixel = 77;
			1662: Pixel = 81;
			1663: Pixel = 112;
			1664: Pixel = 75;
			1665: Pixel = 128;
			1666: Pixel = 160;
			1667: Pixel = 102;
			1668: Pixel = 51;
			1669: Pixel = 55;
			1670: Pixel = 57;
			1671: Pixel = 88;
			1672: Pixel = 119;
			1673: Pixel = 132;
			1674: Pixel = 139;
			1675: Pixel = 139;
			1676: Pixel = 138;
			1677: Pixel = 143;
			1678: Pixel = 145;
			1679: Pixel = 176;
			1680: Pixel = 173;
			1681: Pixel = 143;
			1682: Pixel = 68;
			1683: Pixel = 46;
			1684: Pixel = 75;
			1685: Pixel = 54;
			1686: Pixel = 91;
			1687: Pixel = 137;
			1688: Pixel = 151;
			1689: Pixel = 152;
			1690: Pixel = 148;
			1691: Pixel = 146;
			1692: Pixel = 145;
			1693: Pixel = 133;
			1694: Pixel = 167;
			1695: Pixel = 208;
			1696: Pixel = 208;
			1697: Pixel = 207;
			1698: Pixel = 210;
			1699: Pixel = 212;
			1700: Pixel = 59;
			1701: Pixel = 60;
			1702: Pixel = 97;
			1703: Pixel = 163;
			1704: Pixel = 180;
			1705: Pixel = 169;
			1706: Pixel = 107;
			1707: Pixel = 109;
			1708: Pixel = 94;
			1709: Pixel = 55;
			1710: Pixel = 66;
			1711: Pixel = 101;
			1712: Pixel = 91;
			1713: Pixel = 86;
			1714: Pixel = 118;
			1715: Pixel = 175;
			1716: Pixel = 131;
			1717: Pixel = 64;
			1718: Pixel = 46;
			1719: Pixel = 56;
			1720: Pixel = 60;
			1721: Pixel = 74;
			1722: Pixel = 108;
			1723: Pixel = 126;
			1724: Pixel = 135;
			1725: Pixel = 141;
			1726: Pixel = 116;
			1727: Pixel = 118;
			1728: Pixel = 129;
			1729: Pixel = 141;
			1730: Pixel = 135;
			1731: Pixel = 110;
			1732: Pixel = 43;
			1733: Pixel = 53;
			1734: Pixel = 74;
			1735: Pixel = 59;
			1736: Pixel = 86;
			1737: Pixel = 151;
			1738: Pixel = 152;
			1739: Pixel = 152;
			1740: Pixel = 148;
			1741: Pixel = 146;
			1742: Pixel = 146;
			1743: Pixel = 132;
			1744: Pixel = 177;
			1745: Pixel = 214;
			1746: Pixel = 208;
			1747: Pixel = 211;
			1748: Pixel = 212;
			1749: Pixel = 211;
			1750: Pixel = 53;
			1751: Pixel = 56;
			1752: Pixel = 99;
			1753: Pixel = 159;
			1754: Pixel = 181;
			1755: Pixel = 171;
			1756: Pixel = 98;
			1757: Pixel = 105;
			1758: Pixel = 87;
			1759: Pixel = 60;
			1760: Pixel = 74;
			1761: Pixel = 120;
			1762: Pixel = 96;
			1763: Pixel = 103;
			1764: Pixel = 132;
			1765: Pixel = 165;
			1766: Pixel = 92;
			1767: Pixel = 47;
			1768: Pixel = 52;
			1769: Pixel = 56;
			1770: Pixel = 61;
			1771: Pixel = 66;
			1772: Pixel = 87;
			1773: Pixel = 116;
			1774: Pixel = 127;
			1775: Pixel = 140;
			1776: Pixel = 138;
			1777: Pixel = 126;
			1778: Pixel = 135;
			1779: Pixel = 147;
			1780: Pixel = 146;
			1781: Pixel = 63;
			1782: Pixel = 46;
			1783: Pixel = 54;
			1784: Pixel = 76;
			1785: Pixel = 65;
			1786: Pixel = 88;
			1787: Pixel = 158;
			1788: Pixel = 152;
			1789: Pixel = 154;
			1790: Pixel = 152;
			1791: Pixel = 148;
			1792: Pixel = 144;
			1793: Pixel = 127;
			1794: Pixel = 186;
			1795: Pixel = 218;
			1796: Pixel = 212;
			1797: Pixel = 212;
			1798: Pixel = 206;
			1799: Pixel = 205;
			1800: Pixel = 47;
			1801: Pixel = 59;
			1802: Pixel = 108;
			1803: Pixel = 153;
			1804: Pixel = 179;
			1805: Pixel = 169;
			1806: Pixel = 92;
			1807: Pixel = 89;
			1808: Pixel = 76;
			1809: Pixel = 56;
			1810: Pixel = 69;
			1811: Pixel = 106;
			1812: Pixel = 116;
			1813: Pixel = 108;
			1814: Pixel = 115;
			1815: Pixel = 118;
			1816: Pixel = 45;
			1817: Pixel = 55;
			1818: Pixel = 52;
			1819: Pixel = 51;
			1820: Pixel = 56;
			1821: Pixel = 58;
			1822: Pixel = 64;
			1823: Pixel = 83;
			1824: Pixel = 118;
			1825: Pixel = 135;
			1826: Pixel = 142;
			1827: Pixel = 153;
			1828: Pixel = 160;
			1829: Pixel = 161;
			1830: Pixel = 102;
			1831: Pixel = 44;
			1832: Pixel = 58;
			1833: Pixel = 55;
			1834: Pixel = 82;
			1835: Pixel = 69;
			1836: Pixel = 89;
			1837: Pixel = 161;
			1838: Pixel = 156;
			1839: Pixel = 153;
			1840: Pixel = 152;
			1841: Pixel = 147;
			1842: Pixel = 141;
			1843: Pixel = 123;
			1844: Pixel = 193;
			1845: Pixel = 220;
			1846: Pixel = 212;
			1847: Pixel = 211;
			1848: Pixel = 216;
			1849: Pixel = 215;
			1850: Pixel = 43;
			1851: Pixel = 51;
			1852: Pixel = 104;
			1853: Pixel = 156;
			1854: Pixel = 178;
			1855: Pixel = 165;
			1856: Pixel = 104;
			1857: Pixel = 86;
			1858: Pixel = 67;
			1859: Pixel = 62;
			1860: Pixel = 58;
			1861: Pixel = 101;
			1862: Pixel = 87;
			1863: Pixel = 123;
			1864: Pixel = 132;
			1865: Pixel = 79;
			1866: Pixel = 46;
			1867: Pixel = 61;
			1868: Pixel = 55;
			1869: Pixel = 51;
			1870: Pixel = 51;
			1871: Pixel = 58;
			1872: Pixel = 62;
			1873: Pixel = 60;
			1874: Pixel = 86;
			1875: Pixel = 117;
			1876: Pixel = 136;
			1877: Pixel = 157;
			1878: Pixel = 166;
			1879: Pixel = 159;
			1880: Pixel = 82;
			1881: Pixel = 41;
			1882: Pixel = 55;
			1883: Pixel = 58;
			1884: Pixel = 88;
			1885: Pixel = 75;
			1886: Pixel = 96;
			1887: Pixel = 148;
			1888: Pixel = 133;
			1889: Pixel = 144;
			1890: Pixel = 149;
			1891: Pixel = 148;
			1892: Pixel = 138;
			1893: Pixel = 129;
			1894: Pixel = 206;
			1895: Pixel = 214;
			1896: Pixel = 210;
			1897: Pixel = 211;
			1898: Pixel = 159;
			1899: Pixel = 96;
			1900: Pixel = 65;
			1901: Pixel = 46;
			1902: Pixel = 76;
			1903: Pixel = 150;
			1904: Pixel = 175;
			1905: Pixel = 167;
			1906: Pixel = 121;
			1907: Pixel = 79;
			1908: Pixel = 57;
			1909: Pixel = 63;
			1910: Pixel = 61;
			1911: Pixel = 104;
			1912: Pixel = 98;
			1913: Pixel = 109;
			1914: Pixel = 108;
			1915: Pixel = 126;
			1916: Pixel = 79;
			1917: Pixel = 57;
			1918: Pixel = 57;
			1919: Pixel = 51;
			1920: Pixel = 50;
			1921: Pixel = 56;
			1922: Pixel = 54;
			1923: Pixel = 90;
			1924: Pixel = 124;
			1925: Pixel = 129;
			1926: Pixel = 137;
			1927: Pixel = 146;
			1928: Pixel = 147;
			1929: Pixel = 173;
			1930: Pixel = 185;
			1931: Pixel = 137;
			1932: Pixel = 66;
			1933: Pixel = 43;
			1934: Pixel = 91;
			1935: Pixel = 75;
			1936: Pixel = 103;
			1937: Pixel = 136;
			1938: Pixel = 116;
			1939: Pixel = 115;
			1940: Pixel = 114;
			1941: Pixel = 122;
			1942: Pixel = 118;
			1943: Pixel = 131;
			1944: Pixel = 209;
			1945: Pixel = 207;
			1946: Pixel = 212;
			1947: Pixel = 136;
			1948: Pixel = 46;
			1949: Pixel = 61;
			1950: Pixel = 136;
			1951: Pixel = 95;
			1952: Pixel = 56;
			1953: Pixel = 138;
			1954: Pixel = 175;
			1955: Pixel = 166;
			1956: Pixel = 128;
			1957: Pixel = 58;
			1958: Pixel = 50;
			1959: Pixel = 81;
			1960: Pixel = 80;
			1961: Pixel = 70;
			1962: Pixel = 101;
			1963: Pixel = 86;
			1964: Pixel = 117;
			1965: Pixel = 120;
			1966: Pixel = 96;
			1967: Pixel = 63;
			1968: Pixel = 56;
			1969: Pixel = 53;
			1970: Pixel = 54;
			1971: Pixel = 59;
			1972: Pixel = 59;
			1973: Pixel = 87;
			1974: Pixel = 124;
			1975: Pixel = 129;
			1976: Pixel = 139;
			1977: Pixel = 138;
			1978: Pixel = 150;
			1979: Pixel = 178;
			1980: Pixel = 195;
			1981: Pixel = 210;
			1982: Pixel = 201;
			1983: Pixel = 101;
			1984: Pixel = 65;
			1985: Pixel = 69;
			1986: Pixel = 102;
			1987: Pixel = 151;
			1988: Pixel = 141;
			1989: Pixel = 133;
			1990: Pixel = 119;
			1991: Pixel = 102;
			1992: Pixel = 104;
			1993: Pixel = 120;
			1994: Pixel = 207;
			1995: Pixel = 214;
			1996: Pixel = 138;
			1997: Pixel = 59;
			1998: Pixel = 83;
			1999: Pixel = 92;
			2000: Pixel = 125;
			2001: Pixel = 152;
			2002: Pixel = 72;
			2003: Pixel = 137;
			2004: Pixel = 180;
			2005: Pixel = 170;
			2006: Pixel = 132;
			2007: Pixel = 42;
			2008: Pixel = 57;
			2009: Pixel = 63;
			2010: Pixel = 66;
			2011: Pixel = 60;
			2012: Pixel = 72;
			2013: Pixel = 70;
			2014: Pixel = 111;
			2015: Pixel = 127;
			2016: Pixel = 111;
			2017: Pixel = 80;
			2018: Pixel = 53;
			2019: Pixel = 55;
			2020: Pixel = 56;
			2021: Pixel = 63;
			2022: Pixel = 82;
			2023: Pixel = 82;
			2024: Pixel = 126;
			2025: Pixel = 134;
			2026: Pixel = 139;
			2027: Pixel = 142;
			2028: Pixel = 157;
			2029: Pixel = 169;
			2030: Pixel = 179;
			2031: Pixel = 188;
			2032: Pixel = 207;
			2033: Pixel = 222;
			2034: Pixel = 100;
			2035: Pixel = 46;
			2036: Pixel = 109;
			2037: Pixel = 152;
			2038: Pixel = 143;
			2039: Pixel = 142;
			2040: Pixel = 138;
			2041: Pixel = 129;
			2042: Pixel = 120;
			2043: Pixel = 157;
			2044: Pixel = 221;
			2045: Pixel = 190;
			2046: Pixel = 77;
			2047: Pixel = 91;
			2048: Pixel = 104;
			2049: Pixel = 94;
			2050: Pixel = 71;
			2051: Pixel = 169;
			2052: Pixel = 82;
			2053: Pixel = 133;
			2054: Pixel = 184;
			2055: Pixel = 172;
			2056: Pixel = 111;
			2057: Pixel = 44;
			2058: Pixel = 52;
			2059: Pixel = 52;
			2060: Pixel = 77;
			2061: Pixel = 49;
			2062: Pixel = 67;
			2063: Pixel = 86;
			2064: Pixel = 89;
			2065: Pixel = 132;
			2066: Pixel = 95;
			2067: Pixel = 97;
			2068: Pixel = 52;
			2069: Pixel = 57;
			2070: Pixel = 52;
			2071: Pixel = 61;
			2072: Pixel = 96;
			2073: Pixel = 80;
			2074: Pixel = 131;
			2075: Pixel = 135;
			2076: Pixel = 139;
			2077: Pixel = 144;
			2078: Pixel = 152;
			2079: Pixel = 162;
			2080: Pixel = 174;
			2081: Pixel = 187;
			2082: Pixel = 198;
			2083: Pixel = 218;
			2084: Pixel = 197;
			2085: Pixel = 40;
			2086: Pixel = 111;
			2087: Pixel = 153;
			2088: Pixel = 143;
			2089: Pixel = 140;
			2090: Pixel = 136;
			2091: Pixel = 125;
			2092: Pixel = 147;
			2093: Pixel = 199;
			2094: Pixel = 222;
			2095: Pixel = 145;
			2096: Pixel = 85;
			2097: Pixel = 109;
			2098: Pixel = 96;
			2099: Pixel = 101;
			2100: Pixel = 53;
			2101: Pixel = 165;
			2102: Pixel = 82;
			2103: Pixel = 130;
			2104: Pixel = 185;
			2105: Pixel = 174;
			2106: Pixel = 104;
			2107: Pixel = 46;
			2108: Pixel = 42;
			2109: Pixel = 70;
			2110: Pixel = 76;
			2111: Pixel = 50;
			2112: Pixel = 48;
			2113: Pixel = 70;
			2114: Pixel = 92;
			2115: Pixel = 125;
			2116: Pixel = 125;
			2117: Pixel = 104;
			2118: Pixel = 56;
			2119: Pixel = 58;
			2120: Pixel = 48;
			2121: Pixel = 81;
			2122: Pixel = 109;
			2123: Pixel = 87;
			2124: Pixel = 134;
			2125: Pixel = 136;
			2126: Pixel = 136;
			2127: Pixel = 141;
			2128: Pixel = 148;
			2129: Pixel = 158;
			2130: Pixel = 170;
			2131: Pixel = 184;
			2132: Pixel = 199;
			2133: Pixel = 207;
			2134: Pixel = 228;
			2135: Pixel = 89;
			2136: Pixel = 110;
			2137: Pixel = 154;
			2138: Pixel = 141;
			2139: Pixel = 138;
			2140: Pixel = 129;
			2141: Pixel = 129;
			2142: Pixel = 202;
			2143: Pixel = 217;
			2144: Pixel = 203;
			2145: Pixel = 107;
			2146: Pixel = 99;
			2147: Pixel = 106;
			2148: Pixel = 97;
			2149: Pixel = 99;
			2150: Pixel = 45;
			2151: Pixel = 161;
			2152: Pixel = 94;
			2153: Pixel = 126;
			2154: Pixel = 183;
			2155: Pixel = 172;
			2156: Pixel = 103;
			2157: Pixel = 41;
			2158: Pixel = 50;
			2159: Pixel = 62;
			2160: Pixel = 62;
			2161: Pixel = 51;
			2162: Pixel = 51;
			2163: Pixel = 59;
			2164: Pixel = 88;
			2165: Pixel = 127;
			2166: Pixel = 93;
			2167: Pixel = 76;
			2168: Pixel = 80;
			2169: Pixel = 67;
			2170: Pixel = 50;
			2171: Pixel = 109;
			2172: Pixel = 111;
			2173: Pixel = 95;
			2174: Pixel = 137;
			2175: Pixel = 139;
			2176: Pixel = 136;
			2177: Pixel = 137;
			2178: Pixel = 145;
			2179: Pixel = 154;
			2180: Pixel = 164;
			2181: Pixel = 179;
			2182: Pixel = 195;
			2183: Pixel = 203;
			2184: Pixel = 224;
			2185: Pixel = 147;
			2186: Pixel = 119;
			2187: Pixel = 154;
			2188: Pixel = 139;
			2189: Pixel = 139;
			2190: Pixel = 126;
			2191: Pixel = 139;
			2192: Pixel = 208;
			2193: Pixel = 216;
			2194: Pixel = 166;
			2195: Pixel = 101;
			2196: Pixel = 102;
			2197: Pixel = 96;
			2198: Pixel = 100;
			2199: Pixel = 91;
			2200: Pixel = 40;
			2201: Pixel = 149;
			2202: Pixel = 106;
			2203: Pixel = 125;
			2204: Pixel = 183;
			2205: Pixel = 174;
			2206: Pixel = 112;
			2207: Pixel = 44;
			2208: Pixel = 57;
			2209: Pixel = 52;
			2210: Pixel = 59;
			2211: Pixel = 54;
			2212: Pixel = 54;
			2213: Pixel = 70;
			2214: Pixel = 81;
			2215: Pixel = 92;
			2216: Pixel = 102;
			2217: Pixel = 65;
			2218: Pixel = 51;
			2219: Pixel = 50;
			2220: Pixel = 65;
			2221: Pixel = 124;
			2222: Pixel = 96;
			2223: Pixel = 111;
			2224: Pixel = 143;
			2225: Pixel = 141;
			2226: Pixel = 138;
			2227: Pixel = 136;
			2228: Pixel = 143;
			2229: Pixel = 151;
			2230: Pixel = 159;
			2231: Pixel = 172;
			2232: Pixel = 190;
			2233: Pixel = 202;
			2234: Pixel = 215;
			2235: Pixel = 196;
			2236: Pixel = 124;
			2237: Pixel = 128;
			2238: Pixel = 143;
			2239: Pixel = 146;
			2240: Pixel = 141;
			2241: Pixel = 137;
			2242: Pixel = 165;
			2243: Pixel = 216;
			2244: Pixel = 139;
			2245: Pixel = 95;
			2246: Pixel = 88;
			2247: Pixel = 96;
			2248: Pixel = 95;
			2249: Pixel = 91;
			2250: Pixel = 30;
			2251: Pixel = 143;
			2252: Pixel = 121;
			2253: Pixel = 119;
			2254: Pixel = 181;
			2255: Pixel = 172;
			2256: Pixel = 110;
			2257: Pixel = 49;
			2258: Pixel = 48;
			2259: Pixel = 56;
			2260: Pixel = 61;
			2261: Pixel = 54;
			2262: Pixel = 46;
			2263: Pixel = 73;
			2264: Pixel = 102;
			2265: Pixel = 71;
			2266: Pixel = 81;
			2267: Pixel = 56;
			2268: Pixel = 42;
			2269: Pixel = 44;
			2270: Pixel = 98;
			2271: Pixel = 117;
			2272: Pixel = 80;
			2273: Pixel = 132;
			2274: Pixel = 140;
			2275: Pixel = 142;
			2276: Pixel = 140;
			2277: Pixel = 136;
			2278: Pixel = 140;
			2279: Pixel = 148;
			2280: Pixel = 156;
			2281: Pixel = 166;
			2282: Pixel = 183;
			2283: Pixel = 199;
			2284: Pixel = 209;
			2285: Pixel = 219;
			2286: Pixel = 111;
			2287: Pixel = 76;
			2288: Pixel = 91;
			2289: Pixel = 95;
			2290: Pixel = 123;
			2291: Pixel = 145;
			2292: Pixel = 172;
			2293: Pixel = 205;
			2294: Pixel = 95;
			2295: Pixel = 80;
			2296: Pixel = 92;
			2297: Pixel = 95;
			2298: Pixel = 97;
			2299: Pixel = 72;
			2300: Pixel = 66;
			2301: Pixel = 149;
			2302: Pixel = 141;
			2303: Pixel = 119;
			2304: Pixel = 182;
			2305: Pixel = 173;
			2306: Pixel = 103;
			2307: Pixel = 47;
			2308: Pixel = 50;
			2309: Pixel = 51;
			2310: Pixel = 57;
			2311: Pixel = 56;
			2312: Pixel = 47;
			2313: Pixel = 50;
			2314: Pixel = 94;
			2315: Pixel = 121;
			2316: Pixel = 62;
			2317: Pixel = 40;
			2318: Pixel = 40;
			2319: Pixel = 73;
			2320: Pixel = 117;
			2321: Pixel = 73;
			2322: Pixel = 107;
			2323: Pixel = 140;
			2324: Pixel = 137;
			2325: Pixel = 141;
			2326: Pixel = 142;
			2327: Pixel = 138;
			2328: Pixel = 137;
			2329: Pixel = 142;
			2330: Pixel = 151;
			2331: Pixel = 161;
			2332: Pixel = 175;
			2333: Pixel = 194;
			2334: Pixel = 204;
			2335: Pixel = 221;
			2336: Pixel = 146;
			2337: Pixel = 94;
			2338: Pixel = 91;
			2339: Pixel = 55;
			2340: Pixel = 53;
			2341: Pixel = 176;
			2342: Pixel = 207;
			2343: Pixel = 131;
			2344: Pixel = 55;
			2345: Pixel = 87;
			2346: Pixel = 94;
			2347: Pixel = 88;
			2348: Pixel = 98;
			2349: Pixel = 62;
			2350: Pixel = 91;
			2351: Pixel = 153;
			2352: Pixel = 146;
			2353: Pixel = 122;
			2354: Pixel = 182;
			2355: Pixel = 175;
			2356: Pixel = 94;
			2357: Pixel = 45;
			2358: Pixel = 53;
			2359: Pixel = 51;
			2360: Pixel = 59;
			2361: Pixel = 71;
			2362: Pixel = 58;
			2363: Pixel = 63;
			2364: Pixel = 70;
			2365: Pixel = 102;
			2366: Pixel = 56;
			2367: Pixel = 40;
			2368: Pixel = 47;
			2369: Pixel = 80;
			2370: Pixel = 77;
			2371: Pixel = 97;
			2372: Pixel = 132;
			2373: Pixel = 135;
			2374: Pixel = 139;
			2375: Pixel = 140;
			2376: Pixel = 144;
			2377: Pixel = 142;
			2378: Pixel = 139;
			2379: Pixel = 139;
			2380: Pixel = 146;
			2381: Pixel = 156;
			2382: Pixel = 168;
			2383: Pixel = 185;
			2384: Pixel = 200;
			2385: Pixel = 218;
			2386: Pixel = 179;
			2387: Pixel = 92;
			2388: Pixel = 106;
			2389: Pixel = 90;
			2390: Pixel = 85;
			2391: Pixel = 181;
			2392: Pixel = 131;
			2393: Pixel = 58;
			2394: Pixel = 78;
			2395: Pixel = 97;
			2396: Pixel = 73;
			2397: Pixel = 104;
			2398: Pixel = 91;
			2399: Pixel = 64;
			2400: Pixel = 56;
			2401: Pixel = 131;
			2402: Pixel = 164;
			2403: Pixel = 126;
			2404: Pixel = 181;
			2405: Pixel = 176;
			2406: Pixel = 75;
			2407: Pixel = 44;
			2408: Pixel = 58;
			2409: Pixel = 59;
			2410: Pixel = 59;
			2411: Pixel = 79;
			2412: Pixel = 83;
			2413: Pixel = 65;
			2414: Pixel = 75;
			2415: Pixel = 99;
			2416: Pixel = 52;
			2417: Pixel = 41;
			2418: Pixel = 67;
			2419: Pixel = 92;
			2420: Pixel = 115;
			2421: Pixel = 130;
			2422: Pixel = 128;
			2423: Pixel = 134;
			2424: Pixel = 137;
			2425: Pixel = 140;
			2426: Pixel = 143;
			2427: Pixel = 145;
			2428: Pixel = 144;
			2429: Pixel = 142;
			2430: Pixel = 145;
			2431: Pixel = 153;
			2432: Pixel = 164;
			2433: Pixel = 179;
			2434: Pixel = 192;
			2435: Pixel = 209;
			2436: Pixel = 204;
			2437: Pixel = 95;
			2438: Pixel = 101;
			2439: Pixel = 112;
			2440: Pixel = 115;
			2441: Pixel = 109;
			2442: Pixel = 90;
			2443: Pixel = 86;
			2444: Pixel = 93;
			2445: Pixel = 74;
			2446: Pixel = 90;
			2447: Pixel = 116;
			2448: Pixel = 70;
			2449: Pixel = 53;
			2450: Pixel = 41;
			2451: Pixel = 125;
			2452: Pixel = 197;
			2453: Pixel = 133;
			2454: Pixel = 180;
			2455: Pixel = 170;
			2456: Pixel = 66;
			2457: Pixel = 47;
			2458: Pixel = 62;
			2459: Pixel = 66;
			2460: Pixel = 73;
			2461: Pixel = 72;
			2462: Pixel = 90;
			2463: Pixel = 76;
			2464: Pixel = 63;
			2465: Pixel = 75;
			2466: Pixel = 73;
			2467: Pixel = 60;
			2468: Pixel = 103;
			2469: Pixel = 121;
			2470: Pixel = 125;
			2471: Pixel = 126;
			2472: Pixel = 130;
			2473: Pixel = 133;
			2474: Pixel = 136;
			2475: Pixel = 138;
			2476: Pixel = 142;
			2477: Pixel = 145;
			2478: Pixel = 146;
			2479: Pixel = 148;
			2480: Pixel = 148;
			2481: Pixel = 153;
			2482: Pixel = 162;
			2483: Pixel = 173;
			2484: Pixel = 188;
			2485: Pixel = 200;
			2486: Pixel = 215;
			2487: Pixel = 120;
			2488: Pixel = 90;
			2489: Pixel = 119;
			2490: Pixel = 120;
			2491: Pixel = 119;
			2492: Pixel = 116;
			2493: Pixel = 90;
			2494: Pixel = 82;
			2495: Pixel = 83;
			2496: Pixel = 123;
			2497: Pixel = 86;
			2498: Pixel = 50;
			2499: Pixel = 75;
		endcase
	end
endmodule