module InHandle(
	input wire			nReset,                                                      // Common to all
	input wire			Clk,                                                        // Common to all
	output reg	[7:0]	Pixel,
	output reg			Frame,
	output reg			Line
);

	parameter COLS = 100;
	parameter ROWS = 100;
	
	reg [7:0] col;
	reg [7:0] row;
	
	always @ (posedge Clk or negedge nReset) begin
		if(!nReset) begin   
			Frame <= 0;
	    	Line  <= 0;							
			row <= ROWS-1;
			col <= COLS-1;						// Zero on first pixel	
		end else begin
			if(col == (COLS-1)) begin			// Get ready for next column
	    		Line <= 1;
				col <= 0;
				row <= row + 1;
				if(row == (ROWS-1)) begin		// Get ready for next row
					Frame <= 1;
					row <= 0;
				end
			end else begin
				Line <= 0;
				Frame <= 0;
				col = col + 1;
			end
		end
	end

	always @ (*) begin
		case(col + (row*COLS))


			0: Pixel = 117;
			1: Pixel = 219;
			2: Pixel = 219;
			3: Pixel = 220;
			4: Pixel = 132;
			5: Pixel = 167;
			6: Pixel = 234;
			7: Pixel = 214;
			8: Pixel = 238;
			9: Pixel = 178;
			10: Pixel = 139;
			11: Pixel = 139;
			12: Pixel = 140;
			13: Pixel = 140;
			14: Pixel = 145;
			15: Pixel = 140;
			16: Pixel = 132;
			17: Pixel = 120;
			18: Pixel = 108;
			19: Pixel = 95;
			20: Pixel = 86;
			21: Pixel = 81;
			22: Pixel = 85;
			23: Pixel = 89;
			24: Pixel = 93;
			25: Pixel = 95;
			26: Pixel = 90;
			27: Pixel = 93;
			28: Pixel = 91;
			29: Pixel = 91;
			30: Pixel = 89;
			31: Pixel = 160;
			32: Pixel = 118;
			33: Pixel = 112;
			34: Pixel = 123;
			35: Pixel = 119;
			36: Pixel = 114;
			37: Pixel = 100;
			38: Pixel = 82;
			39: Pixel = 78;
			40: Pixel = 78;
			41: Pixel = 78;
			42: Pixel = 79;
			43: Pixel = 79;
			44: Pixel = 83;
			45: Pixel = 86;
			46: Pixel = 89;
			47: Pixel = 87;
			48: Pixel = 87;
			49: Pixel = 89;
			50: Pixel = 87;
			51: Pixel = 86;
			52: Pixel = 86;
			53: Pixel = 88;
			54: Pixel = 89;
			55: Pixel = 89;
			56: Pixel = 92;
			57: Pixel = 91;
			58: Pixel = 92;
			59: Pixel = 93;
			60: Pixel = 93;
			61: Pixel = 90;
			62: Pixel = 89;
			63: Pixel = 88;
			64: Pixel = 90;
			65: Pixel = 93;
			66: Pixel = 93;
			67: Pixel = 90;
			68: Pixel = 90;
			69: Pixel = 88;
			70: Pixel = 91;
			71: Pixel = 92;
			72: Pixel = 83;
			73: Pixel = 84;
			74: Pixel = 84;
			75: Pixel = 84;
			76: Pixel = 83;
			77: Pixel = 87;
			78: Pixel = 88;
			79: Pixel = 77;
			80: Pixel = 62;
			81: Pixel = 57;
			82: Pixel = 56;
			83: Pixel = 60;
			84: Pixel = 67;
			85: Pixel = 74;
			86: Pixel = 77;
			87: Pixel = 72;
			88: Pixel = 69;
			89: Pixel = 64;
			90: Pixel = 60;
			91: Pixel = 54;
			92: Pixel = 71;
			93: Pixel = 73;
			94: Pixel = 91;
			95: Pixel = 87;
			96: Pixel = 71;
			97: Pixel = 73;
			98: Pixel = 72;
			99: Pixel = 72;
			100: Pixel = 103;
			101: Pixel = 210;
			102: Pixel = 204;
			103: Pixel = 244;
			104: Pixel = 143;
			105: Pixel = 170;
			106: Pixel = 234;
			107: Pixel = 220;
			108: Pixel = 179;
			109: Pixel = 133;
			110: Pixel = 133;
			111: Pixel = 138;
			112: Pixel = 147;
			113: Pixel = 143;
			114: Pixel = 125;
			115: Pixel = 103;
			116: Pixel = 89;
			117: Pixel = 82;
			118: Pixel = 82;
			119: Pixel = 84;
			120: Pixel = 90;
			121: Pixel = 93;
			122: Pixel = 96;
			123: Pixel = 96;
			124: Pixel = 94;
			125: Pixel = 95;
			126: Pixel = 89;
			127: Pixel = 92;
			128: Pixel = 118;
			129: Pixel = 154;
			130: Pixel = 110;
			131: Pixel = 199;
			132: Pixel = 159;
			133: Pixel = 76;
			134: Pixel = 88;
			135: Pixel = 89;
			136: Pixel = 105;
			137: Pixel = 121;
			138: Pixel = 119;
			139: Pixel = 108;
			140: Pixel = 83;
			141: Pixel = 71;
			142: Pixel = 79;
			143: Pixel = 81;
			144: Pixel = 79;
			145: Pixel = 82;
			146: Pixel = 86;
			147: Pixel = 85;
			148: Pixel = 85;
			149: Pixel = 88;
			150: Pixel = 86;
			151: Pixel = 85;
			152: Pixel = 85;
			153: Pixel = 86;
			154: Pixel = 87;
			155: Pixel = 90;
			156: Pixel = 90;
			157: Pixel = 88;
			158: Pixel = 92;
			159: Pixel = 94;
			160: Pixel = 91;
			161: Pixel = 91;
			162: Pixel = 90;
			163: Pixel = 88;
			164: Pixel = 89;
			165: Pixel = 93;
			166: Pixel = 92;
			167: Pixel = 89;
			168: Pixel = 88;
			169: Pixel = 89;
			170: Pixel = 93;
			171: Pixel = 93;
			172: Pixel = 83;
			173: Pixel = 82;
			174: Pixel = 81;
			175: Pixel = 81;
			176: Pixel = 79;
			177: Pixel = 79;
			178: Pixel = 78;
			179: Pixel = 70;
			180: Pixel = 61;
			181: Pixel = 56;
			182: Pixel = 53;
			183: Pixel = 57;
			184: Pixel = 65;
			185: Pixel = 72;
			186: Pixel = 75;
			187: Pixel = 73;
			188: Pixel = 66;
			189: Pixel = 64;
			190: Pixel = 60;
			191: Pixel = 55;
			192: Pixel = 73;
			193: Pixel = 70;
			194: Pixel = 94;
			195: Pixel = 82;
			196: Pixel = 68;
			197: Pixel = 71;
			198: Pixel = 71;
			199: Pixel = 71;
			200: Pixel = 95;
			201: Pixel = 196;
			202: Pixel = 201;
			203: Pixel = 237;
			204: Pixel = 187;
			205: Pixel = 150;
			206: Pixel = 242;
			207: Pixel = 178;
			208: Pixel = 134;
			209: Pixel = 129;
			210: Pixel = 131;
			211: Pixel = 139;
			212: Pixel = 121;
			213: Pixel = 95;
			214: Pixel = 82;
			215: Pixel = 82;
			216: Pixel = 89;
			217: Pixel = 92;
			218: Pixel = 92;
			219: Pixel = 94;
			220: Pixel = 97;
			221: Pixel = 94;
			222: Pixel = 95;
			223: Pixel = 96;
			224: Pixel = 93;
			225: Pixel = 88;
			226: Pixel = 106;
			227: Pixel = 157;
			228: Pixel = 151;
			229: Pixel = 122;
			230: Pixel = 91;
			231: Pixel = 184;
			232: Pixel = 158;
			233: Pixel = 53;
			234: Pixel = 69;
			235: Pixel = 73;
			236: Pixel = 83;
			237: Pixel = 87;
			238: Pixel = 96;
			239: Pixel = 110;
			240: Pixel = 122;
			241: Pixel = 103;
			242: Pixel = 74;
			243: Pixel = 77;
			244: Pixel = 80;
			245: Pixel = 80;
			246: Pixel = 85;
			247: Pixel = 83;
			248: Pixel = 83;
			249: Pixel = 86;
			250: Pixel = 86;
			251: Pixel = 83;
			252: Pixel = 83;
			253: Pixel = 85;
			254: Pixel = 86;
			255: Pixel = 88;
			256: Pixel = 88;
			257: Pixel = 89;
			258: Pixel = 89;
			259: Pixel = 89;
			260: Pixel = 91;
			261: Pixel = 91;
			262: Pixel = 90;
			263: Pixel = 89;
			264: Pixel = 89;
			265: Pixel = 93;
			266: Pixel = 92;
			267: Pixel = 90;
			268: Pixel = 89;
			269: Pixel = 90;
			270: Pixel = 89;
			271: Pixel = 85;
			272: Pixel = 79;
			273: Pixel = 78;
			274: Pixel = 81;
			275: Pixel = 78;
			276: Pixel = 76;
			277: Pixel = 72;
			278: Pixel = 69;
			279: Pixel = 65;
			280: Pixel = 59;
			281: Pixel = 56;
			282: Pixel = 52;
			283: Pixel = 54;
			284: Pixel = 56;
			285: Pixel = 62;
			286: Pixel = 67;
			287: Pixel = 67;
			288: Pixel = 65;
			289: Pixel = 65;
			290: Pixel = 57;
			291: Pixel = 55;
			292: Pixel = 71;
			293: Pixel = 69;
			294: Pixel = 94;
			295: Pixel = 75;
			296: Pixel = 67;
			297: Pixel = 68;
			298: Pixel = 68;
			299: Pixel = 67;
			300: Pixel = 94;
			301: Pixel = 170;
			302: Pixel = 225;
			303: Pixel = 235;
			304: Pixel = 217;
			305: Pixel = 143;
			306: Pixel = 202;
			307: Pixel = 140;
			308: Pixel = 130;
			309: Pixel = 133;
			310: Pixel = 136;
			311: Pixel = 105;
			312: Pixel = 82;
			313: Pixel = 87;
			314: Pixel = 94;
			315: Pixel = 95;
			316: Pixel = 95;
			317: Pixel = 94;
			318: Pixel = 92;
			319: Pixel = 91;
			320: Pixel = 95;
			321: Pixel = 94;
			322: Pixel = 95;
			323: Pixel = 96;
			324: Pixel = 88;
			325: Pixel = 128;
			326: Pixel = 176;
			327: Pixel = 145;
			328: Pixel = 113;
			329: Pixel = 107;
			330: Pixel = 78;
			331: Pixel = 161;
			332: Pixel = 173;
			333: Pixel = 72;
			334: Pixel = 83;
			335: Pixel = 85;
			336: Pixel = 94;
			337: Pixel = 104;
			338: Pixel = 95;
			339: Pixel = 89;
			340: Pixel = 98;
			341: Pixel = 128;
			342: Pixel = 120;
			343: Pixel = 78;
			344: Pixel = 79;
			345: Pixel = 82;
			346: Pixel = 83;
			347: Pixel = 83;
			348: Pixel = 82;
			349: Pixel = 87;
			350: Pixel = 90;
			351: Pixel = 83;
			352: Pixel = 82;
			353: Pixel = 85;
			354: Pixel = 86;
			355: Pixel = 88;
			356: Pixel = 88;
			357: Pixel = 88;
			358: Pixel = 88;
			359: Pixel = 90;
			360: Pixel = 93;
			361: Pixel = 92;
			362: Pixel = 91;
			363: Pixel = 94;
			364: Pixel = 96;
			365: Pixel = 96;
			366: Pixel = 91;
			367: Pixel = 88;
			368: Pixel = 86;
			369: Pixel = 84;
			370: Pixel = 80;
			371: Pixel = 78;
			372: Pixel = 78;
			373: Pixel = 80;
			374: Pixel = 80;
			375: Pixel = 78;
			376: Pixel = 75;
			377: Pixel = 72;
			378: Pixel = 68;
			379: Pixel = 65;
			380: Pixel = 57;
			381: Pixel = 55;
			382: Pixel = 54;
			383: Pixel = 52;
			384: Pixel = 60;
			385: Pixel = 62;
			386: Pixel = 64;
			387: Pixel = 65;
			388: Pixel = 65;
			389: Pixel = 64;
			390: Pixel = 56;
			391: Pixel = 58;
			392: Pixel = 70;
			393: Pixel = 71;
			394: Pixel = 96;
			395: Pixel = 74;
			396: Pixel = 69;
			397: Pixel = 72;
			398: Pixel = 69;
			399: Pixel = 68;
			400: Pixel = 102;
			401: Pixel = 131;
			402: Pixel = 217;
			403: Pixel = 187;
			404: Pixel = 210;
			405: Pixel = 141;
			406: Pixel = 160;
			407: Pixel = 128;
			408: Pixel = 126;
			409: Pixel = 139;
			410: Pixel = 113;
			411: Pixel = 85;
			412: Pixel = 95;
			413: Pixel = 92;
			414: Pixel = 92;
			415: Pixel = 92;
			416: Pixel = 92;
			417: Pixel = 92;
			418: Pixel = 87;
			419: Pixel = 88;
			420: Pixel = 91;
			421: Pixel = 92;
			422: Pixel = 96;
			423: Pixel = 92;
			424: Pixel = 134;
			425: Pixel = 172;
			426: Pixel = 117;
			427: Pixel = 107;
			428: Pixel = 119;
			429: Pixel = 110;
			430: Pixel = 86;
			431: Pixel = 117;
			432: Pixel = 117;
			433: Pixel = 80;
			434: Pixel = 95;
			435: Pixel = 88;
			436: Pixel = 86;
			437: Pixel = 96;
			438: Pixel = 96;
			439: Pixel = 93;
			440: Pixel = 88;
			441: Pixel = 99;
			442: Pixel = 135;
			443: Pixel = 110;
			444: Pixel = 76;
			445: Pixel = 80;
			446: Pixel = 78;
			447: Pixel = 80;
			448: Pixel = 82;
			449: Pixel = 87;
			450: Pixel = 91;
			451: Pixel = 83;
			452: Pixel = 82;
			453: Pixel = 84;
			454: Pixel = 85;
			455: Pixel = 88;
			456: Pixel = 88;
			457: Pixel = 87;
			458: Pixel = 89;
			459: Pixel = 90;
			460: Pixel = 94;
			461: Pixel = 98;
			462: Pixel = 98;
			463: Pixel = 96;
			464: Pixel = 93;
			465: Pixel = 89;
			466: Pixel = 86;
			467: Pixel = 82;
			468: Pixel = 80;
			469: Pixel = 80;
			470: Pixel = 77;
			471: Pixel = 74;
			472: Pixel = 76;
			473: Pixel = 76;
			474: Pixel = 77;
			475: Pixel = 80;
			476: Pixel = 75;
			477: Pixel = 70;
			478: Pixel = 66;
			479: Pixel = 63;
			480: Pixel = 58;
			481: Pixel = 56;
			482: Pixel = 54;
			483: Pixel = 55;
			484: Pixel = 61;
			485: Pixel = 63;
			486: Pixel = 64;
			487: Pixel = 66;
			488: Pixel = 62;
			489: Pixel = 64;
			490: Pixel = 62;
			491: Pixel = 59;
			492: Pixel = 71;
			493: Pixel = 73;
			494: Pixel = 96;
			495: Pixel = 72;
			496: Pixel = 70;
			497: Pixel = 71;
			498: Pixel = 69;
			499: Pixel = 67;
			500: Pixel = 109;
			501: Pixel = 109;
			502: Pixel = 142;
			503: Pixel = 128;
			504: Pixel = 155;
			505: Pixel = 144;
			506: Pixel = 143;
			507: Pixel = 130;
			508: Pixel = 131;
			509: Pixel = 128;
			510: Pixel = 90;
			511: Pixel = 93;
			512: Pixel = 91;
			513: Pixel = 91;
			514: Pixel = 91;
			515: Pixel = 91;
			516: Pixel = 91;
			517: Pixel = 91;
			518: Pixel = 86;
			519: Pixel = 86;
			520: Pixel = 88;
			521: Pixel = 90;
			522: Pixel = 87;
			523: Pixel = 123;
			524: Pixel = 171;
			525: Pixel = 107;
			526: Pixel = 95;
			527: Pixel = 112;
			528: Pixel = 108;
			529: Pixel = 103;
			530: Pixel = 93;
			531: Pixel = 86;
			532: Pixel = 129;
			533: Pixel = 127;
			534: Pixel = 114;
			535: Pixel = 113;
			536: Pixel = 113;
			537: Pixel = 112;
			538: Pixel = 101;
			539: Pixel = 82;
			540: Pixel = 81;
			541: Pixel = 90;
			542: Pixel = 89;
			543: Pixel = 112;
			544: Pixel = 102;
			545: Pixel = 76;
			546: Pixel = 78;
			547: Pixel = 78;
			548: Pixel = 77;
			549: Pixel = 85;
			550: Pixel = 89;
			551: Pixel = 86;
			552: Pixel = 83;
			553: Pixel = 86;
			554: Pixel = 86;
			555: Pixel = 87;
			556: Pixel = 89;
			557: Pixel = 88;
			558: Pixel = 87;
			559: Pixel = 90;
			560: Pixel = 95;
			561: Pixel = 96;
			562: Pixel = 92;
			563: Pixel = 86;
			564: Pixel = 84;
			565: Pixel = 83;
			566: Pixel = 81;
			567: Pixel = 80;
			568: Pixel = 78;
			569: Pixel = 78;
			570: Pixel = 74;
			571: Pixel = 71;
			572: Pixel = 74;
			573: Pixel = 76;
			574: Pixel = 78;
			575: Pixel = 81;
			576: Pixel = 79;
			577: Pixel = 72;
			578: Pixel = 65;
			579: Pixel = 60;
			580: Pixel = 57;
			581: Pixel = 54;
			582: Pixel = 52;
			583: Pixel = 52;
			584: Pixel = 57;
			585: Pixel = 61;
			586: Pixel = 63;
			587: Pixel = 66;
			588: Pixel = 59;
			589: Pixel = 79;
			590: Pixel = 83;
			591: Pixel = 57;
			592: Pixel = 71;
			593: Pixel = 72;
			594: Pixel = 93;
			595: Pixel = 70;
			596: Pixel = 69;
			597: Pixel = 69;
			598: Pixel = 67;
			599: Pixel = 69;
			600: Pixel = 133;
			601: Pixel = 94;
			602: Pixel = 151;
			603: Pixel = 152;
			604: Pixel = 203;
			605: Pixel = 158;
			606: Pixel = 146;
			607: Pixel = 155;
			608: Pixel = 138;
			609: Pixel = 108;
			610: Pixel = 90;
			611: Pixel = 92;
			612: Pixel = 91;
			613: Pixel = 92;
			614: Pixel = 92;
			615: Pixel = 89;
			616: Pixel = 89;
			617: Pixel = 90;
			618: Pixel = 88;
			619: Pixel = 87;
			620: Pixel = 87;
			621: Pixel = 87;
			622: Pixel = 105;
			623: Pixel = 163;
			624: Pixel = 110;
			625: Pixel = 95;
			626: Pixel = 106;
			627: Pixel = 115;
			628: Pixel = 99;
			629: Pixel = 99;
			630: Pixel = 126;
			631: Pixel = 143;
			632: Pixel = 135;
			633: Pixel = 107;
			634: Pixel = 88;
			635: Pixel = 84;
			636: Pixel = 86;
			637: Pixel = 90;
			638: Pixel = 99;
			639: Pixel = 106;
			640: Pixel = 90;
			641: Pixel = 80;
			642: Pixel = 87;
			643: Pixel = 97;
			644: Pixel = 112;
			645: Pixel = 94;
			646: Pixel = 75;
			647: Pixel = 77;
			648: Pixel = 75;
			649: Pixel = 82;
			650: Pixel = 89;
			651: Pixel = 87;
			652: Pixel = 84;
			653: Pixel = 83;
			654: Pixel = 87;
			655: Pixel = 89;
			656: Pixel = 87;
			657: Pixel = 86;
			658: Pixel = 84;
			659: Pixel = 83;
			660: Pixel = 88;
			661: Pixel = 86;
			662: Pixel = 86;
			663: Pixel = 82;
			664: Pixel = 82;
			665: Pixel = 82;
			666: Pixel = 80;
			667: Pixel = 78;
			668: Pixel = 76;
			669: Pixel = 78;
			670: Pixel = 75;
			671: Pixel = 72;
			672: Pixel = 75;
			673: Pixel = 75;
			674: Pixel = 77;
			675: Pixel = 82;
			676: Pixel = 86;
			677: Pixel = 77;
			678: Pixel = 67;
			679: Pixel = 60;
			680: Pixel = 57;
			681: Pixel = 54;
			682: Pixel = 52;
			683: Pixel = 53;
			684: Pixel = 58;
			685: Pixel = 61;
			686: Pixel = 63;
			687: Pixel = 66;
			688: Pixel = 62;
			689: Pixel = 59;
			690: Pixel = 56;
			691: Pixel = 63;
			692: Pixel = 69;
			693: Pixel = 77;
			694: Pixel = 92;
			695: Pixel = 65;
			696: Pixel = 67;
			697: Pixel = 67;
			698: Pixel = 66;
			699: Pixel = 70;
			700: Pixel = 170;
			701: Pixel = 162;
			702: Pixel = 215;
			703: Pixel = 236;
			704: Pixel = 211;
			705: Pixel = 154;
			706: Pixel = 139;
			707: Pixel = 157;
			708: Pixel = 125;
			709: Pixel = 99;
			710: Pixel = 91;
			711: Pixel = 90;
			712: Pixel = 90;
			713: Pixel = 90;
			714: Pixel = 90;
			715: Pixel = 90;
			716: Pixel = 90;
			717: Pixel = 90;
			718: Pixel = 88;
			719: Pixel = 88;
			720: Pixel = 87;
			721: Pixel = 92;
			722: Pixel = 144;
			723: Pixel = 121;
			724: Pixel = 96;
			725: Pixel = 102;
			726: Pixel = 110;
			727: Pixel = 97;
			728: Pixel = 113;
			729: Pixel = 135;
			730: Pixel = 99;
			731: Pixel = 76;
			732: Pixel = 69;
			733: Pixel = 66;
			734: Pixel = 75;
			735: Pixel = 74;
			736: Pixel = 71;
			737: Pixel = 73;
			738: Pixel = 110;
			739: Pixel = 112;
			740: Pixel = 87;
			741: Pixel = 85;
			742: Pixel = 86;
			743: Pixel = 89;
			744: Pixel = 95;
			745: Pixel = 108;
			746: Pixel = 82;
			747: Pixel = 76;
			748: Pixel = 74;
			749: Pixel = 79;
			750: Pixel = 89;
			751: Pixel = 88;
			752: Pixel = 85;
			753: Pixel = 88;
			754: Pixel = 89;
			755: Pixel = 89;
			756: Pixel = 87;
			757: Pixel = 86;
			758: Pixel = 82;
			759: Pixel = 81;
			760: Pixel = 83;
			761: Pixel = 85;
			762: Pixel = 84;
			763: Pixel = 81;
			764: Pixel = 81;
			765: Pixel = 82;
			766: Pixel = 80;
			767: Pixel = 77;
			768: Pixel = 75;
			769: Pixel = 76;
			770: Pixel = 76;
			771: Pixel = 74;
			772: Pixel = 75;
			773: Pixel = 74;
			774: Pixel = 75;
			775: Pixel = 82;
			776: Pixel = 85;
			777: Pixel = 78;
			778: Pixel = 70;
			779: Pixel = 62;
			780: Pixel = 59;
			781: Pixel = 57;
			782: Pixel = 54;
			783: Pixel = 54;
			784: Pixel = 59;
			785: Pixel = 61;
			786: Pixel = 64;
			787: Pixel = 67;
			788: Pixel = 66;
			789: Pixel = 63;
			790: Pixel = 55;
			791: Pixel = 64;
			792: Pixel = 68;
			793: Pixel = 82;
			794: Pixel = 92;
			795: Pixel = 65;
			796: Pixel = 69;
			797: Pixel = 69;
			798: Pixel = 67;
			799: Pixel = 68;
			800: Pixel = 173;
			801: Pixel = 255;
			802: Pixel = 212;
			803: Pixel = 221;
			804: Pixel = 201;
			805: Pixel = 128;
			806: Pixel = 110;
			807: Pixel = 95;
			808: Pixel = 113;
			809: Pixel = 94;
			810: Pixel = 91;
			811: Pixel = 88;
			812: Pixel = 88;
			813: Pixel = 88;
			814: Pixel = 89;
			815: Pixel = 89;
			816: Pixel = 91;
			817: Pixel = 89;
			818: Pixel = 87;
			819: Pixel = 87;
			820: Pixel = 83;
			821: Pixel = 121;
			822: Pixel = 164;
			823: Pixel = 108;
			824: Pixel = 101;
			825: Pixel = 94;
			826: Pixel = 89;
			827: Pixel = 107;
			828: Pixel = 117;
			829: Pixel = 75;
			830: Pixel = 63;
			831: Pixel = 73;
			832: Pixel = 71;
			833: Pixel = 67;
			834: Pixel = 73;
			835: Pixel = 74;
			836: Pixel = 68;
			837: Pixel = 77;
			838: Pixel = 98;
			839: Pixel = 111;
			840: Pixel = 103;
			841: Pixel = 75;
			842: Pixel = 78;
			843: Pixel = 82;
			844: Pixel = 83;
			845: Pixel = 101;
			846: Pixel = 99;
			847: Pixel = 74;
			848: Pixel = 73;
			849: Pixel = 77;
			850: Pixel = 89;
			851: Pixel = 90;
			852: Pixel = 89;
			853: Pixel = 89;
			854: Pixel = 85;
			855: Pixel = 86;
			856: Pixel = 84;
			857: Pixel = 83;
			858: Pixel = 81;
			859: Pixel = 79;
			860: Pixel = 81;
			861: Pixel = 81;
			862: Pixel = 82;
			863: Pixel = 82;
			864: Pixel = 82;
			865: Pixel = 82;
			866: Pixel = 80;
			867: Pixel = 77;
			868: Pixel = 76;
			869: Pixel = 77;
			870: Pixel = 76;
			871: Pixel = 72;
			872: Pixel = 70;
			873: Pixel = 70;
			874: Pixel = 76;
			875: Pixel = 79;
			876: Pixel = 74;
			877: Pixel = 71;
			878: Pixel = 69;
			879: Pixel = 61;
			880: Pixel = 54;
			881: Pixel = 55;
			882: Pixel = 53;
			883: Pixel = 55;
			884: Pixel = 55;
			885: Pixel = 59;
			886: Pixel = 64;
			887: Pixel = 66;
			888: Pixel = 68;
			889: Pixel = 65;
			890: Pixel = 56;
			891: Pixel = 64;
			892: Pixel = 67;
			893: Pixel = 84;
			894: Pixel = 87;
			895: Pixel = 64;
			896: Pixel = 70;
			897: Pixel = 71;
			898: Pixel = 68;
			899: Pixel = 66;
			900: Pixel = 168;
			901: Pixel = 197;
			902: Pixel = 158;
			903: Pixel = 136;
			904: Pixel = 155;
			905: Pixel = 129;
			906: Pixel = 115;
			907: Pixel = 120;
			908: Pixel = 115;
			909: Pixel = 88;
			910: Pixel = 90;
			911: Pixel = 88;
			912: Pixel = 87;
			913: Pixel = 87;
			914: Pixel = 89;
			915: Pixel = 89;
			916: Pixel = 88;
			917: Pixel = 86;
			918: Pixel = 86;
			919: Pixel = 84;
			920: Pixel = 95;
			921: Pixel = 134;
			922: Pixel = 116;
			923: Pixel = 105;
			924: Pixel = 95;
			925: Pixel = 88;
			926: Pixel = 121;
			927: Pixel = 146;
			928: Pixel = 88;
			929: Pixel = 71;
			930: Pixel = 70;
			931: Pixel = 72;
			932: Pixel = 69;
			933: Pixel = 65;
			934: Pixel = 71;
			935: Pixel = 72;
			936: Pixel = 67;
			937: Pixel = 78;
			938: Pixel = 83;
			939: Pixel = 115;
			940: Pixel = 119;
			941: Pixel = 73;
			942: Pixel = 61;
			943: Pixel = 70;
			944: Pixel = 80;
			945: Pixel = 88;
			946: Pixel = 104;
			947: Pixel = 85;
			948: Pixel = 74;
			949: Pixel = 78;
			950: Pixel = 84;
			951: Pixel = 88;
			952: Pixel = 86;
			953: Pixel = 87;
			954: Pixel = 83;
			955: Pixel = 83;
			956: Pixel = 82;
			957: Pixel = 81;
			958: Pixel = 80;
			959: Pixel = 79;
			960: Pixel = 81;
			961: Pixel = 84;
			962: Pixel = 82;
			963: Pixel = 83;
			964: Pixel = 83;
			965: Pixel = 81;
			966: Pixel = 78;
			967: Pixel = 75;
			968: Pixel = 75;
			969: Pixel = 79;
			970: Pixel = 77;
			971: Pixel = 72;
			972: Pixel = 70;
			973: Pixel = 73;
			974: Pixel = 76;
			975: Pixel = 70;
			976: Pixel = 66;
			977: Pixel = 65;
			978: Pixel = 64;
			979: Pixel = 59;
			980: Pixel = 54;
			981: Pixel = 54;
			982: Pixel = 54;
			983: Pixel = 54;
			984: Pixel = 56;
			985: Pixel = 59;
			986: Pixel = 64;
			987: Pixel = 65;
			988: Pixel = 63;
			989: Pixel = 64;
			990: Pixel = 55;
			991: Pixel = 67;
			992: Pixel = 68;
			993: Pixel = 89;
			994: Pixel = 83;
			995: Pixel = 65;
			996: Pixel = 73;
			997: Pixel = 72;
			998: Pixel = 68;
			999: Pixel = 64;
			1000: Pixel = 134;
			1001: Pixel = 148;
			1002: Pixel = 155;
			1003: Pixel = 141;
			1004: Pixel = 158;
			1005: Pixel = 140;
			1006: Pixel = 107;
			1007: Pixel = 121;
			1008: Pixel = 118;
			1009: Pixel = 86;
			1010: Pixel = 88;
			1011: Pixel = 88;
			1012: Pixel = 86;
			1013: Pixel = 88;
			1014: Pixel = 87;
			1015: Pixel = 88;
			1016: Pixel = 86;
			1017: Pixel = 84;
			1018: Pixel = 84;
			1019: Pixel = 81;
			1020: Pixel = 123;
			1021: Pixel = 116;
			1022: Pixel = 88;
			1023: Pixel = 92;
			1024: Pixel = 83;
			1025: Pixel = 103;
			1026: Pixel = 155;
			1027: Pixel = 137;
			1028: Pixel = 113;
			1029: Pixel = 88;
			1030: Pixel = 66;
			1031: Pixel = 70;
			1032: Pixel = 70;
			1033: Pixel = 64;
			1034: Pixel = 65;
			1035: Pixel = 69;
			1036: Pixel = 69;
			1037: Pixel = 65;
			1038: Pixel = 67;
			1039: Pixel = 88;
			1040: Pixel = 137;
			1041: Pixel = 68;
			1042: Pixel = 61;
			1043: Pixel = 61;
			1044: Pixel = 69;
			1045: Pixel = 85;
			1046: Pixel = 97;
			1047: Pixel = 99;
			1048: Pixel = 72;
			1049: Pixel = 76;
			1050: Pixel = 79;
			1051: Pixel = 85;
			1052: Pixel = 83;
			1053: Pixel = 84;
			1054: Pixel = 83;
			1055: Pixel = 81;
			1056: Pixel = 81;
			1057: Pixel = 80;
			1058: Pixel = 80;
			1059: Pixel = 79;
			1060: Pixel = 80;
			1061: Pixel = 84;
			1062: Pixel = 81;
			1063: Pixel = 82;
			1064: Pixel = 82;
			1065: Pixel = 80;
			1066: Pixel = 78;
			1067: Pixel = 74;
			1068: Pixel = 75;
			1069: Pixel = 76;
			1070: Pixel = 78;
			1071: Pixel = 76;
			1072: Pixel = 72;
			1073: Pixel = 75;
			1074: Pixel = 69;
			1075: Pixel = 62;
			1076: Pixel = 60;
			1077: Pixel = 61;
			1078: Pixel = 61;
			1079: Pixel = 56;
			1080: Pixel = 54;
			1081: Pixel = 54;
			1082: Pixel = 54;
			1083: Pixel = 53;
			1084: Pixel = 56;
			1085: Pixel = 56;
			1086: Pixel = 62;
			1087: Pixel = 64;
			1088: Pixel = 62;
			1089: Pixel = 61;
			1090: Pixel = 54;
			1091: Pixel = 67;
			1092: Pixel = 66;
			1093: Pixel = 93;
			1094: Pixel = 78;
			1095: Pixel = 64;
			1096: Pixel = 72;
			1097: Pixel = 72;
			1098: Pixel = 70;
			1099: Pixel = 64;
			1100: Pixel = 151;
			1101: Pixel = 194;
			1102: Pixel = 165;
			1103: Pixel = 121;
			1104: Pixel = 101;
			1105: Pixel = 108;
			1106: Pixel = 109;
			1107: Pixel = 110;
			1108: Pixel = 119;
			1109: Pixel = 89;
			1110: Pixel = 87;
			1111: Pixel = 88;
			1112: Pixel = 88;
			1113: Pixel = 90;
			1114: Pixel = 88;
			1115: Pixel = 88;
			1116: Pixel = 86;
			1117: Pixel = 84;
			1118: Pixel = 82;
			1119: Pixel = 90;
			1120: Pixel = 131;
			1121: Pixel = 97;
			1122: Pixel = 95;
			1123: Pixel = 84;
			1124: Pixel = 91;
			1125: Pixel = 113;
			1126: Pixel = 88;
			1127: Pixel = 144;
			1128: Pixel = 137;
			1129: Pixel = 92;
			1130: Pixel = 70;
			1131: Pixel = 70;
			1132: Pixel = 72;
			1133: Pixel = 74;
			1134: Pixel = 90;
			1135: Pixel = 99;
			1136: Pixel = 95;
			1137: Pixel = 69;
			1138: Pixel = 59;
			1139: Pixel = 72;
			1140: Pixel = 74;
			1141: Pixel = 65;
			1142: Pixel = 61;
			1143: Pixel = 62;
			1144: Pixel = 61;
			1145: Pixel = 76;
			1146: Pixel = 94;
			1147: Pixel = 108;
			1148: Pixel = 82;
			1149: Pixel = 72;
			1150: Pixel = 79;
			1151: Pixel = 85;
			1152: Pixel = 85;
			1153: Pixel = 83;
			1154: Pixel = 83;
			1155: Pixel = 80;
			1156: Pixel = 82;
			1157: Pixel = 83;
			1158: Pixel = 82;
			1159: Pixel = 80;
			1160: Pixel = 79;
			1161: Pixel = 80;
			1162: Pixel = 81;
			1163: Pixel = 81;
			1164: Pixel = 83;
			1165: Pixel = 81;
			1166: Pixel = 78;
			1167: Pixel = 75;
			1168: Pixel = 74;
			1169: Pixel = 74;
			1170: Pixel = 76;
			1171: Pixel = 78;
			1172: Pixel = 75;
			1173: Pixel = 69;
			1174: Pixel = 64;
			1175: Pixel = 62;
			1176: Pixel = 61;
			1177: Pixel = 58;
			1178: Pixel = 58;
			1179: Pixel = 54;
			1180: Pixel = 55;
			1181: Pixel = 56;
			1182: Pixel = 55;
			1183: Pixel = 54;
			1184: Pixel = 56;
			1185: Pixel = 58;
			1186: Pixel = 62;
			1187: Pixel = 65;
			1188: Pixel = 63;
			1189: Pixel = 61;
			1190: Pixel = 58;
			1191: Pixel = 69;
			1192: Pixel = 70;
			1193: Pixel = 97;
			1194: Pixel = 77;
			1195: Pixel = 69;
			1196: Pixel = 76;
			1197: Pixel = 74;
			1198: Pixel = 76;
			1199: Pixel = 61;
			1200: Pixel = 130;
			1201: Pixel = 140;
			1202: Pixel = 147;
			1203: Pixel = 112;
			1204: Pixel = 64;
			1205: Pixel = 94;
			1206: Pixel = 113;
			1207: Pixel = 107;
			1208: Pixel = 118;
			1209: Pixel = 92;
			1210: Pixel = 87;
			1211: Pixel = 88;
			1212: Pixel = 87;
			1213: Pixel = 89;
			1214: Pixel = 88;
			1215: Pixel = 86;
			1216: Pixel = 86;
			1217: Pixel = 84;
			1218: Pixel = 77;
			1219: Pixel = 109;
			1220: Pixel = 118;
			1221: Pixel = 95;
			1222: Pixel = 89;
			1223: Pixel = 82;
			1224: Pixel = 101;
			1225: Pixel = 78;
			1226: Pixel = 83;
			1227: Pixel = 126;
			1228: Pixel = 145;
			1229: Pixel = 87;
			1230: Pixel = 64;
			1231: Pixel = 77;
			1232: Pixel = 127;
			1233: Pixel = 168;
			1234: Pixel = 185;
			1235: Pixel = 177;
			1236: Pixel = 162;
			1237: Pixel = 105;
			1238: Pixel = 61;
			1239: Pixel = 62;
			1240: Pixel = 61;
			1241: Pixel = 61;
			1242: Pixel = 61;
			1243: Pixel = 61;
			1244: Pixel = 61;
			1245: Pixel = 63;
			1246: Pixel = 87;
			1247: Pixel = 112;
			1248: Pixel = 94;
			1249: Pixel = 69;
			1250: Pixel = 77;
			1251: Pixel = 84;
			1252: Pixel = 83;
			1253: Pixel = 83;
			1254: Pixel = 84;
			1255: Pixel = 81;
			1256: Pixel = 84;
			1257: Pixel = 84;
			1258: Pixel = 81;
			1259: Pixel = 79;
			1260: Pixel = 80;
			1261: Pixel = 81;
			1262: Pixel = 83;
			1263: Pixel = 82;
			1264: Pixel = 85;
			1265: Pixel = 78;
			1266: Pixel = 78;
			1267: Pixel = 75;
			1268: Pixel = 75;
			1269: Pixel = 74;
			1270: Pixel = 73;
			1271: Pixel = 73;
			1272: Pixel = 71;
			1273: Pixel = 65;
			1274: Pixel = 62;
			1275: Pixel = 60;
			1276: Pixel = 58;
			1277: Pixel = 57;
			1278: Pixel = 56;
			1279: Pixel = 52;
			1280: Pixel = 53;
			1281: Pixel = 55;
			1282: Pixel = 55;
			1283: Pixel = 55;
			1284: Pixel = 57;
			1285: Pixel = 62;
			1286: Pixel = 61;
			1287: Pixel = 63;
			1288: Pixel = 66;
			1289: Pixel = 62;
			1290: Pixel = 59;
			1291: Pixel = 70;
			1292: Pixel = 72;
			1293: Pixel = 97;
			1294: Pixel = 73;
			1295: Pixel = 71;
			1296: Pixel = 76;
			1297: Pixel = 82;
			1298: Pixel = 81;
			1299: Pixel = 57;
			1300: Pixel = 79;
			1301: Pixel = 108;
			1302: Pixel = 137;
			1303: Pixel = 109;
			1304: Pixel = 71;
			1305: Pixel = 87;
			1306: Pixel = 113;
			1307: Pixel = 103;
			1308: Pixel = 117;
			1309: Pixel = 95;
			1310: Pixel = 85;
			1311: Pixel = 88;
			1312: Pixel = 86;
			1313: Pixel = 86;
			1314: Pixel = 86;
			1315: Pixel = 85;
			1316: Pixel = 82;
			1317: Pixel = 80;
			1318: Pixel = 80;
			1319: Pixel = 117;
			1320: Pixel = 103;
			1321: Pixel = 92;
			1322: Pixel = 79;
			1323: Pixel = 91;
			1324: Pixel = 86;
			1325: Pixel = 63;
			1326: Pixel = 72;
			1327: Pixel = 91;
			1328: Pixel = 182;
			1329: Pixel = 101;
			1330: Pixel = 74;
			1331: Pixel = 152;
			1332: Pixel = 207;
			1333: Pixel = 214;
			1334: Pixel = 206;
			1335: Pixel = 188;
			1336: Pixel = 168;
			1337: Pixel = 117;
			1338: Pixel = 72;
			1339: Pixel = 60;
			1340: Pixel = 67;
			1341: Pixel = 59;
			1342: Pixel = 60;
			1343: Pixel = 60;
			1344: Pixel = 60;
			1345: Pixel = 61;
			1346: Pixel = 72;
			1347: Pixel = 106;
			1348: Pixel = 105;
			1349: Pixel = 71;
			1350: Pixel = 76;
			1351: Pixel = 83;
			1352: Pixel = 82;
			1353: Pixel = 85;
			1354: Pixel = 84;
			1355: Pixel = 81;
			1356: Pixel = 82;
			1357: Pixel = 82;
			1358: Pixel = 82;
			1359: Pixel = 81;
			1360: Pixel = 79;
			1361: Pixel = 79;
			1362: Pixel = 81;
			1363: Pixel = 79;
			1364: Pixel = 80;
			1365: Pixel = 76;
			1366: Pixel = 79;
			1367: Pixel = 77;
			1368: Pixel = 73;
			1369: Pixel = 71;
			1370: Pixel = 69;
			1371: Pixel = 70;
			1372: Pixel = 66;
			1373: Pixel = 63;
			1374: Pixel = 60;
			1375: Pixel = 58;
			1376: Pixel = 56;
			1377: Pixel = 55;
			1378: Pixel = 53;
			1379: Pixel = 54;
			1380: Pixel = 52;
			1381: Pixel = 53;
			1382: Pixel = 54;
			1383: Pixel = 55;
			1384: Pixel = 59;
			1385: Pixel = 63;
			1386: Pixel = 62;
			1387: Pixel = 61;
			1388: Pixel = 65;
			1389: Pixel = 60;
			1390: Pixel = 60;
			1391: Pixel = 68;
			1392: Pixel = 72;
			1393: Pixel = 98;
			1394: Pixel = 72;
			1395: Pixel = 74;
			1396: Pixel = 81;
			1397: Pixel = 87;
			1398: Pixel = 75;
			1399: Pixel = 53;
			1400: Pixel = 79;
			1401: Pixel = 98;
			1402: Pixel = 115;
			1403: Pixel = 129;
			1404: Pixel = 72;
			1405: Pixel = 78;
			1406: Pixel = 113;
			1407: Pixel = 102;
			1408: Pixel = 111;
			1409: Pixel = 99;
			1410: Pixel = 83;
			1411: Pixel = 87;
			1412: Pixel = 85;
			1413: Pixel = 85;
			1414: Pixel = 84;
			1415: Pixel = 83;
			1416: Pixel = 80;
			1417: Pixel = 77;
			1418: Pixel = 90;
			1419: Pixel = 119;
			1420: Pixel = 94;
			1421: Pixel = 85;
			1422: Pixel = 77;
			1423: Pixel = 98;
			1424: Pixel = 66;
			1425: Pixel = 64;
			1426: Pixel = 60;
			1427: Pixel = 71;
			1428: Pixel = 83;
			1429: Pixel = 77;
			1430: Pixel = 102;
			1431: Pixel = 194;
			1432: Pixel = 193;
			1433: Pixel = 202;
			1434: Pixel = 227;
			1435: Pixel = 222;
			1436: Pixel = 210;
			1437: Pixel = 141;
			1438: Pixel = 91;
			1439: Pixel = 85;
			1440: Pixel = 84;
			1441: Pixel = 67;
			1442: Pixel = 59;
			1443: Pixel = 60;
			1444: Pixel = 61;
			1445: Pixel = 62;
			1446: Pixel = 65;
			1447: Pixel = 77;
			1448: Pixel = 113;
			1449: Pixel = 81;
			1450: Pixel = 73;
			1451: Pixel = 83;
			1452: Pixel = 84;
			1453: Pixel = 86;
			1454: Pixel = 84;
			1455: Pixel = 83;
			1456: Pixel = 83;
			1457: Pixel = 83;
			1458: Pixel = 83;
			1459: Pixel = 82;
			1460: Pixel = 82;
			1461: Pixel = 82;
			1462: Pixel = 81;
			1463: Pixel = 80;
			1464: Pixel = 79;
			1465: Pixel = 78;
			1466: Pixel = 78;
			1467: Pixel = 76;
			1468: Pixel = 74;
			1469: Pixel = 71;
			1470: Pixel = 69;
			1471: Pixel = 68;
			1472: Pixel = 64;
			1473: Pixel = 64;
			1474: Pixel = 61;
			1475: Pixel = 58;
			1476: Pixel = 56;
			1477: Pixel = 54;
			1478: Pixel = 54;
			1479: Pixel = 53;
			1480: Pixel = 53;
			1481: Pixel = 56;
			1482: Pixel = 55;
			1483: Pixel = 59;
			1484: Pixel = 63;
			1485: Pixel = 64;
			1486: Pixel = 65;
			1487: Pixel = 61;
			1488: Pixel = 64;
			1489: Pixel = 61;
			1490: Pixel = 63;
			1491: Pixel = 69;
			1492: Pixel = 76;
			1493: Pixel = 92;
			1494: Pixel = 73;
			1495: Pixel = 82;
			1496: Pixel = 87;
			1497: Pixel = 80;
			1498: Pixel = 71;
			1499: Pixel = 53;
			1500: Pixel = 80;
			1501: Pixel = 151;
			1502: Pixel = 117;
			1503: Pixel = 117;
			1504: Pixel = 64;
			1505: Pixel = 71;
			1506: Pixel = 109;
			1507: Pixel = 105;
			1508: Pixel = 108;
			1509: Pixel = 103;
			1510: Pixel = 82;
			1511: Pixel = 84;
			1512: Pixel = 85;
			1513: Pixel = 85;
			1514: Pixel = 86;
			1515: Pixel = 84;
			1516: Pixel = 83;
			1517: Pixel = 78;
			1518: Pixel = 103;
			1519: Pixel = 114;
			1520: Pixel = 95;
			1521: Pixel = 79;
			1522: Pixel = 85;
			1523: Pixel = 85;
			1524: Pixel = 59;
			1525: Pixel = 64;
			1526: Pixel = 62;
			1527: Pixel = 59;
			1528: Pixel = 59;
			1529: Pixel = 58;
			1530: Pixel = 99;
			1531: Pixel = 182;
			1532: Pixel = 230;
			1533: Pixel = 248;
			1534: Pixel = 251;
			1535: Pixel = 238;
			1536: Pixel = 228;
			1537: Pixel = 173;
			1538: Pixel = 109;
			1539: Pixel = 110;
			1540: Pixel = 88;
			1541: Pixel = 78;
			1542: Pixel = 64;
			1543: Pixel = 59;
			1544: Pixel = 61;
			1545: Pixel = 63;
			1546: Pixel = 62;
			1547: Pixel = 76;
			1548: Pixel = 118;
			1549: Pixel = 91;
			1550: Pixel = 72;
			1551: Pixel = 81;
			1552: Pixel = 85;
			1553: Pixel = 94;
			1554: Pixel = 83;
			1555: Pixel = 86;
			1556: Pixel = 88;
			1557: Pixel = 85;
			1558: Pixel = 84;
			1559: Pixel = 83;
			1560: Pixel = 83;
			1561: Pixel = 81;
			1562: Pixel = 81;
			1563: Pixel = 82;
			1564: Pixel = 81;
			1565: Pixel = 78;
			1566: Pixel = 78;
			1567: Pixel = 76;
			1568: Pixel = 76;
			1569: Pixel = 73;
			1570: Pixel = 72;
			1571: Pixel = 70;
			1572: Pixel = 67;
			1573: Pixel = 65;
			1574: Pixel = 62;
			1575: Pixel = 57;
			1576: Pixel = 56;
			1577: Pixel = 53;
			1578: Pixel = 53;
			1579: Pixel = 55;
			1580: Pixel = 56;
			1581: Pixel = 58;
			1582: Pixel = 61;
			1583: Pixel = 65;
			1584: Pixel = 66;
			1585: Pixel = 66;
			1586: Pixel = 67;
			1587: Pixel = 66;
			1588: Pixel = 67;
			1589: Pixel = 62;
			1590: Pixel = 65;
			1591: Pixel = 70;
			1592: Pixel = 81;
			1593: Pixel = 96;
			1594: Pixel = 79;
			1595: Pixel = 93;
			1596: Pixel = 88;
			1597: Pixel = 75;
			1598: Pixel = 71;
			1599: Pixel = 52;
			1600: Pixel = 116;
			1601: Pixel = 158;
			1602: Pixel = 129;
			1603: Pixel = 105;
			1604: Pixel = 74;
			1605: Pixel = 61;
			1606: Pixel = 102;
			1607: Pixel = 107;
			1608: Pixel = 108;
			1609: Pixel = 109;
			1610: Pixel = 82;
			1611: Pixel = 85;
			1612: Pixel = 85;
			1613: Pixel = 86;
			1614: Pixel = 85;
			1615: Pixel = 84;
			1616: Pixel = 82;
			1617: Pixel = 79;
			1618: Pixel = 110;
			1619: Pixel = 109;
			1620: Pixel = 93;
			1621: Pixel = 72;
			1622: Pixel = 85;
			1623: Pixel = 70;
			1624: Pixel = 61;
			1625: Pixel = 61;
			1626: Pixel = 61;
			1627: Pixel = 60;
			1628: Pixel = 71;
			1629: Pixel = 81;
			1630: Pixel = 120;
			1631: Pixel = 213;
			1632: Pixel = 254;
			1633: Pixel = 235;
			1634: Pixel = 215;
			1635: Pixel = 194;
			1636: Pixel = 168;
			1637: Pixel = 139;
			1638: Pixel = 123;
			1639: Pixel = 127;
			1640: Pixel = 99;
			1641: Pixel = 87;
			1642: Pixel = 72;
			1643: Pixel = 60;
			1644: Pixel = 61;
			1645: Pixel = 62;
			1646: Pixel = 64;
			1647: Pixel = 69;
			1648: Pixel = 108;
			1649: Pixel = 98;
			1650: Pixel = 74;
			1651: Pixel = 76;
			1652: Pixel = 144;
			1653: Pixel = 208;
			1654: Pixel = 126;
			1655: Pixel = 82;
			1656: Pixel = 88;
			1657: Pixel = 85;
			1658: Pixel = 85;
			1659: Pixel = 85;
			1660: Pixel = 81;
			1661: Pixel = 81;
			1662: Pixel = 80;
			1663: Pixel = 80;
			1664: Pixel = 80;
			1665: Pixel = 78;
			1666: Pixel = 78;
			1667: Pixel = 77;
			1668: Pixel = 77;
			1669: Pixel = 73;
			1670: Pixel = 73;
			1671: Pixel = 71;
			1672: Pixel = 70;
			1673: Pixel = 69;
			1674: Pixel = 63;
			1675: Pixel = 60;
			1676: Pixel = 56;
			1677: Pixel = 55;
			1678: Pixel = 53;
			1679: Pixel = 56;
			1680: Pixel = 58;
			1681: Pixel = 61;
			1682: Pixel = 67;
			1683: Pixel = 67;
			1684: Pixel = 67;
			1685: Pixel = 66;
			1686: Pixel = 66;
			1687: Pixel = 65;
			1688: Pixel = 64;
			1689: Pixel = 61;
			1690: Pixel = 66;
			1691: Pixel = 70;
			1692: Pixel = 85;
			1693: Pixel = 97;
			1694: Pixel = 94;
			1695: Pixel = 100;
			1696: Pixel = 86;
			1697: Pixel = 75;
			1698: Pixel = 71;
			1699: Pixel = 58;
			1700: Pixel = 186;
			1701: Pixel = 115;
			1702: Pixel = 117;
			1703: Pixel = 126;
			1704: Pixel = 113;
			1705: Pixel = 65;
			1706: Pixel = 92;
			1707: Pixel = 109;
			1708: Pixel = 106;
			1709: Pixel = 116;
			1710: Pixel = 84;
			1711: Pixel = 84;
			1712: Pixel = 86;
			1713: Pixel = 84;
			1714: Pixel = 83;
			1715: Pixel = 82;
			1716: Pixel = 80;
			1717: Pixel = 80;
			1718: Pixel = 111;
			1719: Pixel = 103;
			1720: Pixel = 86;
			1721: Pixel = 68;
			1722: Pixel = 79;
			1723: Pixel = 61;
			1724: Pixel = 62;
			1725: Pixel = 61;
			1726: Pixel = 57;
			1727: Pixel = 72;
			1728: Pixel = 114;
			1729: Pixel = 123;
			1730: Pixel = 155;
			1731: Pixel = 220;
			1732: Pixel = 227;
			1733: Pixel = 190;
			1734: Pixel = 193;
			1735: Pixel = 178;
			1736: Pixel = 151;
			1737: Pixel = 120;
			1738: Pixel = 110;
			1739: Pixel = 103;
			1740: Pixel = 96;
			1741: Pixel = 88;
			1742: Pixel = 78;
			1743: Pixel = 61;
			1744: Pixel = 58;
			1745: Pixel = 60;
			1746: Pixel = 59;
			1747: Pixel = 63;
			1748: Pixel = 97;
			1749: Pixel = 102;
			1750: Pixel = 69;
			1751: Pixel = 100;
			1752: Pixel = 220;
			1753: Pixel = 236;
			1754: Pixel = 222;
			1755: Pixel = 132;
			1756: Pixel = 92;
			1757: Pixel = 87;
			1758: Pixel = 86;
			1759: Pixel = 85;
			1760: Pixel = 81;
			1761: Pixel = 80;
			1762: Pixel = 81;
			1763: Pixel = 80;
			1764: Pixel = 81;
			1765: Pixel = 77;
			1766: Pixel = 76;
			1767: Pixel = 76;
			1768: Pixel = 77;
			1769: Pixel = 73;
			1770: Pixel = 74;
			1771: Pixel = 70;
			1772: Pixel = 71;
			1773: Pixel = 69;
			1774: Pixel = 66;
			1775: Pixel = 61;
			1776: Pixel = 55;
			1777: Pixel = 54;
			1778: Pixel = 55;
			1779: Pixel = 55;
			1780: Pixel = 57;
			1781: Pixel = 65;
			1782: Pixel = 67;
			1783: Pixel = 66;
			1784: Pixel = 68;
			1785: Pixel = 67;
			1786: Pixel = 66;
			1787: Pixel = 62;
			1788: Pixel = 61;
			1789: Pixel = 58;
			1790: Pixel = 67;
			1791: Pixel = 69;
			1792: Pixel = 89;
			1793: Pixel = 100;
			1794: Pixel = 95;
			1795: Pixel = 89;
			1796: Pixel = 81;
			1797: Pixel = 72;
			1798: Pixel = 67;
			1799: Pixel = 57;
			1800: Pixel = 173;
			1801: Pixel = 105;
			1802: Pixel = 156;
			1803: Pixel = 158;
			1804: Pixel = 101;
			1805: Pixel = 54;
			1806: Pixel = 81;
			1807: Pixel = 112;
			1808: Pixel = 103;
			1809: Pixel = 116;
			1810: Pixel = 89;
			1811: Pixel = 82;
			1812: Pixel = 85;
			1813: Pixel = 84;
			1814: Pixel = 83;
			1815: Pixel = 82;
			1816: Pixel = 78;
			1817: Pixel = 80;
			1818: Pixel = 112;
			1819: Pixel = 99;
			1820: Pixel = 81;
			1821: Pixel = 69;
			1822: Pixel = 72;
			1823: Pixel = 59;
			1824: Pixel = 61;
			1825: Pixel = 59;
			1826: Pixel = 58;
			1827: Pixel = 98;
			1828: Pixel = 136;
			1829: Pixel = 171;
			1830: Pixel = 231;
			1831: Pixel = 203;
			1832: Pixel = 172;
			1833: Pixel = 180;
			1834: Pixel = 183;
			1835: Pixel = 165;
			1836: Pixel = 140;
			1837: Pixel = 114;
			1838: Pixel = 106;
			1839: Pixel = 97;
			1840: Pixel = 82;
			1841: Pixel = 81;
			1842: Pixel = 79;
			1843: Pixel = 64;
			1844: Pixel = 61;
			1845: Pixel = 65;
			1846: Pixel = 82;
			1847: Pixel = 69;
			1848: Pixel = 87;
			1849: Pixel = 102;
			1850: Pixel = 65;
			1851: Pixel = 152;
			1852: Pixel = 231;
			1853: Pixel = 219;
			1854: Pixel = 230;
			1855: Pixel = 214;
			1856: Pixel = 140;
			1857: Pixel = 106;
			1858: Pixel = 91;
			1859: Pixel = 84;
			1860: Pixel = 83;
			1861: Pixel = 80;
			1862: Pixel = 80;
			1863: Pixel = 82;
			1864: Pixel = 80;
			1865: Pixel = 78;
			1866: Pixel = 77;
			1867: Pixel = 77;
			1868: Pixel = 78;
			1869: Pixel = 80;
			1870: Pixel = 77;
			1871: Pixel = 70;
			1872: Pixel = 71;
			1873: Pixel = 72;
			1874: Pixel = 68;
			1875: Pixel = 62;
			1876: Pixel = 57;
			1877: Pixel = 56;
			1878: Pixel = 56;
			1879: Pixel = 56;
			1880: Pixel = 58;
			1881: Pixel = 66;
			1882: Pixel = 68;
			1883: Pixel = 70;
			1884: Pixel = 65;
			1885: Pixel = 68;
			1886: Pixel = 66;
			1887: Pixel = 62;
			1888: Pixel = 65;
			1889: Pixel = 65;
			1890: Pixel = 68;
			1891: Pixel = 71;
			1892: Pixel = 95;
			1893: Pixel = 99;
			1894: Pixel = 83;
			1895: Pixel = 81;
			1896: Pixel = 76;
			1897: Pixel = 73;
			1898: Pixel = 66;
			1899: Pixel = 57;
			1900: Pixel = 160;
			1901: Pixel = 167;
			1902: Pixel = 190;
			1903: Pixel = 184;
			1904: Pixel = 149;
			1905: Pixel = 119;
			1906: Pixel = 80;
			1907: Pixel = 108;
			1908: Pixel = 104;
			1909: Pixel = 115;
			1910: Pixel = 96;
			1911: Pixel = 81;
			1912: Pixel = 83;
			1913: Pixel = 84;
			1914: Pixel = 83;
			1915: Pixel = 82;
			1916: Pixel = 79;
			1917: Pixel = 82;
			1918: Pixel = 118;
			1919: Pixel = 105;
			1920: Pixel = 80;
			1921: Pixel = 71;
			1922: Pixel = 66;
			1923: Pixel = 60;
			1924: Pixel = 60;
			1925: Pixel = 56;
			1926: Pixel = 65;
			1927: Pixel = 114;
			1928: Pixel = 145;
			1929: Pixel = 194;
			1930: Pixel = 214;
			1931: Pixel = 159;
			1932: Pixel = 138;
			1933: Pixel = 155;
			1934: Pixel = 162;
			1935: Pixel = 158;
			1936: Pixel = 145;
			1937: Pixel = 118;
			1938: Pixel = 110;
			1939: Pixel = 103;
			1940: Pixel = 81;
			1941: Pixel = 73;
			1942: Pixel = 74;
			1943: Pixel = 71;
			1944: Pixel = 61;
			1945: Pixel = 123;
			1946: Pixel = 127;
			1947: Pixel = 79;
			1948: Pixel = 84;
			1949: Pixel = 100;
			1950: Pixel = 77;
			1951: Pixel = 192;
			1952: Pixel = 222;
			1953: Pixel = 222;
			1954: Pixel = 221;
			1955: Pixel = 225;
			1956: Pixel = 217;
			1957: Pixel = 147;
			1958: Pixel = 110;
			1959: Pixel = 89;
			1960: Pixel = 84;
			1961: Pixel = 81;
			1962: Pixel = 81;
			1963: Pixel = 82;
			1964: Pixel = 82;
			1965: Pixel = 81;
			1966: Pixel = 80;
			1967: Pixel = 79;
			1968: Pixel = 80;
			1969: Pixel = 85;
			1970: Pixel = 80;
			1971: Pixel = 74;
			1972: Pixel = 71;
			1973: Pixel = 67;
			1974: Pixel = 73;
			1975: Pixel = 68;
			1976: Pixel = 62;
			1977: Pixel = 59;
			1978: Pixel = 57;
			1979: Pixel = 56;
			1980: Pixel = 61;
			1981: Pixel = 69;
			1982: Pixel = 71;
			1983: Pixel = 74;
			1984: Pixel = 82;
			1985: Pixel = 65;
			1986: Pixel = 71;
			1987: Pixel = 57;
			1988: Pixel = 107;
			1989: Pixel = 98;
			1990: Pixel = 65;
			1991: Pixel = 73;
			1992: Pixel = 98;
			1993: Pixel = 92;
			1994: Pixel = 78;
			1995: Pixel = 82;
			1996: Pixel = 77;
			1997: Pixel = 81;
			1998: Pixel = 66;
			1999: Pixel = 57;
			2000: Pixel = 189;
			2001: Pixel = 147;
			2002: Pixel = 144;
			2003: Pixel = 139;
			2004: Pixel = 121;
			2005: Pixel = 136;
			2006: Pixel = 154;
			2007: Pixel = 121;
			2008: Pixel = 106;
			2009: Pixel = 117;
			2010: Pixel = 105;
			2011: Pixel = 82;
			2012: Pixel = 85;
			2013: Pixel = 85;
			2014: Pixel = 83;
			2015: Pixel = 81;
			2016: Pixel = 79;
			2017: Pixel = 83;
			2018: Pixel = 129;
			2019: Pixel = 118;
			2020: Pixel = 75;
			2021: Pixel = 71;
			2022: Pixel = 62;
			2023: Pixel = 61;
			2024: Pixel = 60;
			2025: Pixel = 59;
			2026: Pixel = 72;
			2027: Pixel = 119;
			2028: Pixel = 150;
			2029: Pixel = 202;
			2030: Pixel = 173;
			2031: Pixel = 133;
			2032: Pixel = 120;
			2033: Pixel = 132;
			2034: Pixel = 162;
			2035: Pixel = 165;
			2036: Pixel = 154;
			2037: Pixel = 132;
			2038: Pixel = 117;
			2039: Pixel = 114;
			2040: Pixel = 92;
			2041: Pixel = 73;
			2042: Pixel = 68;
			2043: Pixel = 74;
			2044: Pixel = 70;
			2045: Pixel = 111;
			2046: Pixel = 112;
			2047: Pixel = 100;
			2048: Pixel = 84;
			2049: Pixel = 95;
			2050: Pixel = 108;
			2051: Pixel = 212;
			2052: Pixel = 212;
			2053: Pixel = 220;
			2054: Pixel = 222;
			2055: Pixel = 221;
			2056: Pixel = 233;
			2057: Pixel = 223;
			2058: Pixel = 143;
			2059: Pixel = 107;
			2060: Pixel = 86;
			2061: Pixel = 85;
			2062: Pixel = 83;
			2063: Pixel = 81;
			2064: Pixel = 84;
			2065: Pixel = 84;
			2066: Pixel = 83;
			2067: Pixel = 83;
			2068: Pixel = 82;
			2069: Pixel = 80;
			2070: Pixel = 76;
			2071: Pixel = 73;
			2072: Pixel = 65;
			2073: Pixel = 51;
			2074: Pixel = 69;
			2075: Pixel = 67;
			2076: Pixel = 62;
			2077: Pixel = 62;
			2078: Pixel = 61;
			2079: Pixel = 57;
			2080: Pixel = 62;
			2081: Pixel = 69;
			2082: Pixel = 71;
			2083: Pixel = 70;
			2084: Pixel = 100;
			2085: Pixel = 63;
			2086: Pixel = 64;
			2087: Pixel = 56;
			2088: Pixel = 70;
			2089: Pixel = 72;
			2090: Pixel = 72;
			2091: Pixel = 74;
			2092: Pixel = 97;
			2093: Pixel = 89;
			2094: Pixel = 76;
			2095: Pixel = 82;
			2096: Pixel = 81;
			2097: Pixel = 85;
			2098: Pixel = 64;
			2099: Pixel = 59;
			2100: Pixel = 219;
			2101: Pixel = 177;
			2102: Pixel = 127;
			2103: Pixel = 115;
			2104: Pixel = 110;
			2105: Pixel = 149;
			2106: Pixel = 241;
			2107: Pixel = 142;
			2108: Pixel = 102;
			2109: Pixel = 117;
			2110: Pixel = 114;
			2111: Pixel = 80;
			2112: Pixel = 83;
			2113: Pixel = 84;
			2114: Pixel = 83;
			2115: Pixel = 79;
			2116: Pixel = 78;
			2117: Pixel = 86;
			2118: Pixel = 114;
			2119: Pixel = 97;
			2120: Pixel = 76;
			2121: Pixel = 67;
			2122: Pixel = 60;
			2123: Pixel = 59;
			2124: Pixel = 57;
			2125: Pixel = 58;
			2126: Pixel = 78;
			2127: Pixel = 115;
			2128: Pixel = 141;
			2129: Pixel = 165;
			2130: Pixel = 131;
			2131: Pixel = 126;
			2132: Pixel = 123;
			2133: Pixel = 121;
			2134: Pixel = 151;
			2135: Pixel = 168;
			2136: Pixel = 162;
			2137: Pixel = 153;
			2138: Pixel = 138;
			2139: Pixel = 128;
			2140: Pixel = 106;
			2141: Pixel = 79;
			2142: Pixel = 64;
			2143: Pixel = 60;
			2144: Pixel = 53;
			2145: Pixel = 67;
			2146: Pixel = 114;
			2147: Pixel = 121;
			2148: Pixel = 87;
			2149: Pixel = 88;
			2150: Pixel = 154;
			2151: Pixel = 216;
			2152: Pixel = 212;
			2153: Pixel = 216;
			2154: Pixel = 218;
			2155: Pixel = 221;
			2156: Pixel = 222;
			2157: Pixel = 244;
			2158: Pixel = 215;
			2159: Pixel = 160;
			2160: Pixel = 112;
			2161: Pixel = 84;
			2162: Pixel = 85;
			2163: Pixel = 87;
			2164: Pixel = 87;
			2165: Pixel = 85;
			2166: Pixel = 82;
			2167: Pixel = 79;
			2168: Pixel = 77;
			2169: Pixel = 74;
			2170: Pixel = 76;
			2171: Pixel = 67;
			2172: Pixel = 45;
			2173: Pixel = 29;
			2174: Pixel = 48;
			2175: Pixel = 68;
			2176: Pixel = 75;
			2177: Pixel = 83;
			2178: Pixel = 62;
			2179: Pixel = 59;
			2180: Pixel = 64;
			2181: Pixel = 70;
			2182: Pixel = 75;
			2183: Pixel = 75;
			2184: Pixel = 63;
			2185: Pixel = 64;
			2186: Pixel = 57;
			2187: Pixel = 50;
			2188: Pixel = 64;
			2189: Pixel = 61;
			2190: Pixel = 71;
			2191: Pixel = 78;
			2192: Pixel = 99;
			2193: Pixel = 85;
			2194: Pixel = 77;
			2195: Pixel = 83;
			2196: Pixel = 85;
			2197: Pixel = 86;
			2198: Pixel = 58;
			2199: Pixel = 78;
			2200: Pixel = 231;
			2201: Pixel = 175;
			2202: Pixel = 104;
			2203: Pixel = 132;
			2204: Pixel = 166;
			2205: Pixel = 196;
			2206: Pixel = 236;
			2207: Pixel = 157;
			2208: Pixel = 106;
			2209: Pixel = 117;
			2210: Pixel = 124;
			2211: Pixel = 84;
			2212: Pixel = 81;
			2213: Pixel = 84;
			2214: Pixel = 84;
			2215: Pixel = 78;
			2216: Pixel = 79;
			2217: Pixel = 84;
			2218: Pixel = 112;
			2219: Pixel = 99;
			2220: Pixel = 76;
			2221: Pixel = 62;
			2222: Pixel = 59;
			2223: Pixel = 59;
			2224: Pixel = 57;
			2225: Pixel = 60;
			2226: Pixel = 79;
			2227: Pixel = 106;
			2228: Pixel = 122;
			2229: Pixel = 128;
			2230: Pixel = 109;
			2231: Pixel = 119;
			2232: Pixel = 131;
			2233: Pixel = 122;
			2234: Pixel = 152;
			2235: Pixel = 176;
			2236: Pixel = 173;
			2237: Pixel = 168;
			2238: Pixel = 160;
			2239: Pixel = 149;
			2240: Pixel = 129;
			2241: Pixel = 93;
			2242: Pixel = 60;
			2243: Pixel = 54;
			2244: Pixel = 52;
			2245: Pixel = 56;
			2246: Pixel = 83;
			2247: Pixel = 128;
			2248: Pixel = 77;
			2249: Pixel = 114;
			2250: Pixel = 214;
			2251: Pixel = 205;
			2252: Pixel = 171;
			2253: Pixel = 218;
			2254: Pixel = 219;
			2255: Pixel = 218;
			2256: Pixel = 223;
			2257: Pixel = 236;
			2258: Pixel = 249;
			2259: Pixel = 232;
			2260: Pixel = 193;
			2261: Pixel = 128;
			2262: Pixel = 84;
			2263: Pixel = 82;
			2264: Pixel = 79;
			2265: Pixel = 78;
			2266: Pixel = 76;
			2267: Pixel = 76;
			2268: Pixel = 75;
			2269: Pixel = 74;
			2270: Pixel = 76;
			2271: Pixel = 58;
			2272: Pixel = 52;
			2273: Pixel = 79;
			2274: Pixel = 44;
			2275: Pixel = 53;
			2276: Pixel = 91;
			2277: Pixel = 95;
			2278: Pixel = 60;
			2279: Pixel = 70;
			2280: Pixel = 72;
			2281: Pixel = 78;
			2282: Pixel = 80;
			2283: Pixel = 80;
			2284: Pixel = 77;
			2285: Pixel = 72;
			2286: Pixel = 70;
			2287: Pixel = 57;
			2288: Pixel = 69;
			2289: Pixel = 64;
			2290: Pixel = 70;
			2291: Pixel = 78;
			2292: Pixel = 102;
			2293: Pixel = 87;
			2294: Pixel = 80;
			2295: Pixel = 85;
			2296: Pixel = 87;
			2297: Pixel = 77;
			2298: Pixel = 59;
			2299: Pixel = 114;
			2300: Pixel = 214;
			2301: Pixel = 160;
			2302: Pixel = 113;
			2303: Pixel = 187;
			2304: Pixel = 214;
			2305: Pixel = 224;
			2306: Pixel = 236;
			2307: Pixel = 209;
			2308: Pixel = 111;
			2309: Pixel = 113;
			2310: Pixel = 132;
			2311: Pixel = 93;
			2312: Pixel = 81;
			2313: Pixel = 85;
			2314: Pixel = 81;
			2315: Pixel = 76;
			2316: Pixel = 78;
			2317: Pixel = 81;
			2318: Pixel = 110;
			2319: Pixel = 100;
			2320: Pixel = 78;
			2321: Pixel = 61;
			2322: Pixel = 58;
			2323: Pixel = 56;
			2324: Pixel = 57;
			2325: Pixel = 62;
			2326: Pixel = 73;
			2327: Pixel = 96;
			2328: Pixel = 110;
			2329: Pixel = 110;
			2330: Pixel = 99;
			2331: Pixel = 114;
			2332: Pixel = 129;
			2333: Pixel = 142;
			2334: Pixel = 173;
			2335: Pixel = 188;
			2336: Pixel = 188;
			2337: Pixel = 178;
			2338: Pixel = 173;
			2339: Pixel = 167;
			2340: Pixel = 149;
			2341: Pixel = 118;
			2342: Pixel = 76;
			2343: Pixel = 61;
			2344: Pixel = 61;
			2345: Pixel = 60;
			2346: Pixel = 70;
			2347: Pixel = 63;
			2348: Pixel = 98;
			2349: Pixel = 212;
			2350: Pixel = 248;
			2351: Pixel = 178;
			2352: Pixel = 67;
			2353: Pixel = 179;
			2354: Pixel = 225;
			2355: Pixel = 217;
			2356: Pixel = 219;
			2357: Pixel = 237;
			2358: Pixel = 244;
			2359: Pixel = 245;
			2360: Pixel = 245;
			2361: Pixel = 219;
			2362: Pixel = 98;
			2363: Pixel = 76;
			2364: Pixel = 79;
			2365: Pixel = 77;
			2366: Pixel = 76;
			2367: Pixel = 77;
			2368: Pixel = 74;
			2369: Pixel = 73;
			2370: Pixel = 74;
			2371: Pixel = 53;
			2372: Pixel = 60;
			2373: Pixel = 105;
			2374: Pixel = 102;
			2375: Pixel = 54;
			2376: Pixel = 64;
			2377: Pixel = 70;
			2378: Pixel = 72;
			2379: Pixel = 77;
			2380: Pixel = 73;
			2381: Pixel = 70;
			2382: Pixel = 77;
			2383: Pixel = 73;
			2384: Pixel = 75;
			2385: Pixel = 75;
			2386: Pixel = 72;
			2387: Pixel = 56;
			2388: Pixel = 72;
			2389: Pixel = 64;
			2390: Pixel = 67;
			2391: Pixel = 73;
			2392: Pixel = 98;
			2393: Pixel = 88;
			2394: Pixel = 85;
			2395: Pixel = 90;
			2396: Pixel = 91;
			2397: Pixel = 54;
			2398: Pixel = 59;
			2399: Pixel = 90;
			2400: Pixel = 161;
			2401: Pixel = 184;
			2402: Pixel = 125;
			2403: Pixel = 176;
			2404: Pixel = 181;
			2405: Pixel = 189;
			2406: Pixel = 238;
			2407: Pixel = 230;
			2408: Pixel = 128;
			2409: Pixel = 109;
			2410: Pixel = 133;
			2411: Pixel = 101;
			2412: Pixel = 81;
			2413: Pixel = 86;
			2414: Pixel = 82;
			2415: Pixel = 79;
			2416: Pixel = 77;
			2417: Pixel = 81;
			2418: Pixel = 109;
			2419: Pixel = 102;
			2420: Pixel = 81;
			2421: Pixel = 59;
			2422: Pixel = 57;
			2423: Pixel = 65;
			2424: Pixel = 67;
			2425: Pixel = 67;
			2426: Pixel = 69;
			2427: Pixel = 86;
			2428: Pixel = 101;
			2429: Pixel = 93;
			2430: Pixel = 91;
			2431: Pixel = 106;
			2432: Pixel = 121;
			2433: Pixel = 155;
			2434: Pixel = 193;
			2435: Pixel = 204;
			2436: Pixel = 199;
			2437: Pixel = 190;
			2438: Pixel = 180;
			2439: Pixel = 177;
			2440: Pixel = 162;
			2441: Pixel = 139;
			2442: Pixel = 108;
			2443: Pixel = 65;
			2444: Pixel = 65;
			2445: Pixel = 70;
			2446: Pixel = 68;
			2447: Pixel = 76;
			2448: Pixel = 217;
			2449: Pixel = 236;
			2450: Pixel = 238;
			2451: Pixel = 196;
			2452: Pixel = 97;
			2453: Pixel = 90;
			2454: Pixel = 220;
			2455: Pixel = 223;
			2456: Pixel = 221;
			2457: Pixel = 229;
			2458: Pixel = 207;
			2459: Pixel = 223;
			2460: Pixel = 237;
			2461: Pixel = 252;
			2462: Pixel = 123;
			2463: Pixel = 71;
			2464: Pixel = 82;
			2465: Pixel = 79;
			2466: Pixel = 79;
			2467: Pixel = 77;
			2468: Pixel = 74;
			2469: Pixel = 74;
			2470: Pixel = 70;
			2471: Pixel = 49;
			2472: Pixel = 36;
			2473: Pixel = 102;
			2474: Pixel = 152;
			2475: Pixel = 85;
			2476: Pixel = 66;
			2477: Pixel = 72;
			2478: Pixel = 69;
			2479: Pixel = 67;
			2480: Pixel = 70;
			2481: Pixel = 73;
			2482: Pixel = 77;
			2483: Pixel = 75;
			2484: Pixel = 77;
			2485: Pixel = 78;
			2486: Pixel = 73;
			2487: Pixel = 59;
			2488: Pixel = 77;
			2489: Pixel = 69;
			2490: Pixel = 67;
			2491: Pixel = 70;
			2492: Pixel = 95;
			2493: Pixel = 94;
			2494: Pixel = 90;
			2495: Pixel = 92;
			2496: Pixel = 93;
			2497: Pixel = 59;
			2498: Pixel = 51;
			2499: Pixel = 64;
			2500: Pixel = 144;
			2501: Pixel = 135;
			2502: Pixel = 139;
			2503: Pixel = 137;
			2504: Pixel = 87;
			2505: Pixel = 145;
			2506: Pixel = 244;
			2507: Pixel = 237;
			2508: Pixel = 149;
			2509: Pixel = 106;
			2510: Pixel = 130;
			2511: Pixel = 111;
			2512: Pixel = 79;
			2513: Pixel = 83;
			2514: Pixel = 82;
			2515: Pixel = 76;
			2516: Pixel = 75;
			2517: Pixel = 78;
			2518: Pixel = 106;
			2519: Pixel = 103;
			2520: Pixel = 82;
			2521: Pixel = 56;
			2522: Pixel = 71;
			2523: Pixel = 109;
			2524: Pixel = 93;
			2525: Pixel = 71;
			2526: Pixel = 71;
			2527: Pixel = 80;
			2528: Pixel = 91;
			2529: Pixel = 82;
			2530: Pixel = 84;
			2531: Pixel = 98;
			2532: Pixel = 118;
			2533: Pixel = 161;
			2534: Pixel = 202;
			2535: Pixel = 222;
			2536: Pixel = 210;
			2537: Pixel = 198;
			2538: Pixel = 184;
			2539: Pixel = 181;
			2540: Pixel = 175;
			2541: Pixel = 151;
			2542: Pixel = 129;
			2543: Pixel = 85;
			2544: Pixel = 65;
			2545: Pixel = 73;
			2546: Pixel = 57;
			2547: Pixel = 140;
			2548: Pixel = 252;
			2549: Pixel = 218;
			2550: Pixel = 231;
			2551: Pixel = 226;
			2552: Pixel = 145;
			2553: Pixel = 120;
			2554: Pixel = 228;
			2555: Pixel = 223;
			2556: Pixel = 228;
			2557: Pixel = 197;
			2558: Pixel = 155;
			2559: Pixel = 180;
			2560: Pixel = 195;
			2561: Pixel = 221;
			2562: Pixel = 111;
			2563: Pixel = 72;
			2564: Pixel = 81;
			2565: Pixel = 77;
			2566: Pixel = 77;
			2567: Pixel = 76;
			2568: Pixel = 73;
			2569: Pixel = 70;
			2570: Pixel = 66;
			2571: Pixel = 59;
			2572: Pixel = 22;
			2573: Pixel = 80;
			2574: Pixel = 163;
			2575: Pixel = 114;
			2576: Pixel = 65;
			2577: Pixel = 71;
			2578: Pixel = 64;
			2579: Pixel = 66;
			2580: Pixel = 68;
			2581: Pixel = 74;
			2582: Pixel = 77;
			2583: Pixel = 76;
			2584: Pixel = 78;
			2585: Pixel = 78;
			2586: Pixel = 73;
			2587: Pixel = 63;
			2588: Pixel = 80;
			2589: Pixel = 70;
			2590: Pixel = 66;
			2591: Pixel = 68;
			2592: Pixel = 91;
			2593: Pixel = 98;
			2594: Pixel = 93;
			2595: Pixel = 95;
			2596: Pixel = 98;
			2597: Pixel = 79;
			2598: Pixel = 48;
			2599: Pixel = 53;
			2600: Pixel = 208;
			2601: Pixel = 93;
			2602: Pixel = 123;
			2603: Pixel = 151;
			2604: Pixel = 87;
			2605: Pixel = 153;
			2606: Pixel = 245;
			2607: Pixel = 242;
			2608: Pixel = 176;
			2609: Pixel = 108;
			2610: Pixel = 130;
			2611: Pixel = 122;
			2612: Pixel = 81;
			2613: Pixel = 84;
			2614: Pixel = 83;
			2615: Pixel = 77;
			2616: Pixel = 76;
			2617: Pixel = 74;
			2618: Pixel = 99;
			2619: Pixel = 106;
			2620: Pixel = 85;
			2621: Pixel = 58;
			2622: Pixel = 86;
			2623: Pixel = 117;
			2624: Pixel = 117;
			2625: Pixel = 73;
			2626: Pixel = 55;
			2627: Pixel = 68;
			2628: Pixel = 79;
			2629: Pixel = 74;
			2630: Pixel = 75;
			2631: Pixel = 93;
			2632: Pixel = 118;
			2633: Pixel = 161;
			2634: Pixel = 202;
			2635: Pixel = 232;
			2636: Pixel = 228;
			2637: Pixel = 205;
			2638: Pixel = 192;
			2639: Pixel = 185;
			2640: Pixel = 188;
			2641: Pixel = 201;
			2642: Pixel = 164;
			2643: Pixel = 116;
			2644: Pixel = 73;
			2645: Pixel = 85;
			2646: Pixel = 155;
			2647: Pixel = 220;
			2648: Pixel = 223;
			2649: Pixel = 218;
			2650: Pixel = 211;
			2651: Pixel = 193;
			2652: Pixel = 164;
			2653: Pixel = 200;
			2654: Pixel = 245;
			2655: Pixel = 232;
			2656: Pixel = 225;
			2657: Pixel = 170;
			2658: Pixel = 144;
			2659: Pixel = 146;
			2660: Pixel = 156;
			2661: Pixel = 171;
			2662: Pixel = 89;
			2663: Pixel = 77;
			2664: Pixel = 80;
			2665: Pixel = 78;
			2666: Pixel = 77;
			2667: Pixel = 76;
			2668: Pixel = 73;
			2669: Pixel = 70;
			2670: Pixel = 67;
			2671: Pixel = 76;
			2672: Pixel = 51;
			2673: Pixel = 67;
			2674: Pixel = 153;
			2675: Pixel = 137;
			2676: Pixel = 75;
			2677: Pixel = 69;
			2678: Pixel = 64;
			2679: Pixel = 64;
			2680: Pixel = 66;
			2681: Pixel = 70;
			2682: Pixel = 77;
			2683: Pixel = 79;
			2684: Pixel = 79;
			2685: Pixel = 79;
			2686: Pixel = 75;
			2687: Pixel = 64;
			2688: Pixel = 82;
			2689: Pixel = 75;
			2690: Pixel = 65;
			2691: Pixel = 66;
			2692: Pixel = 92;
			2693: Pixel = 103;
			2694: Pixel = 96;
			2695: Pixel = 98;
			2696: Pixel = 101;
			2697: Pixel = 81;
			2698: Pixel = 49;
			2699: Pixel = 49;
			2700: Pixel = 171;
			2701: Pixel = 122;
			2702: Pixel = 119;
			2703: Pixel = 178;
			2704: Pixel = 181;
			2705: Pixel = 214;
			2706: Pixel = 236;
			2707: Pixel = 239;
			2708: Pixel = 198;
			2709: Pixel = 113;
			2710: Pixel = 130;
			2711: Pixel = 132;
			2712: Pixel = 87;
			2713: Pixel = 86;
			2714: Pixel = 85;
			2715: Pixel = 80;
			2716: Pixel = 78;
			2717: Pixel = 75;
			2718: Pixel = 92;
			2719: Pixel = 109;
			2720: Pixel = 89;
			2721: Pixel = 62;
			2722: Pixel = 63;
			2723: Pixel = 123;
			2724: Pixel = 137;
			2725: Pixel = 83;
			2726: Pixel = 48;
			2727: Pixel = 62;
			2728: Pixel = 76;
			2729: Pixel = 69;
			2730: Pixel = 68;
			2731: Pixel = 84;
			2732: Pixel = 117;
			2733: Pixel = 152;
			2734: Pixel = 193;
			2735: Pixel = 228;
			2736: Pixel = 240;
			2737: Pixel = 219;
			2738: Pixel = 201;
			2739: Pixel = 191;
			2740: Pixel = 213;
			2741: Pixel = 255;
			2742: Pixel = 182;
			2743: Pixel = 130;
			2744: Pixel = 130;
			2745: Pixel = 205;
			2746: Pixel = 242;
			2747: Pixel = 230;
			2748: Pixel = 223;
			2749: Pixel = 225;
			2750: Pixel = 227;
			2751: Pixel = 232;
			2752: Pixel = 227;
			2753: Pixel = 208;
			2754: Pixel = 234;
			2755: Pixel = 250;
			2756: Pixel = 220;
			2757: Pixel = 157;
			2758: Pixel = 147;
			2759: Pixel = 141;
			2760: Pixel = 142;
			2761: Pixel = 123;
			2762: Pixel = 80;
			2763: Pixel = 80;
			2764: Pixel = 79;
			2765: Pixel = 77;
			2766: Pixel = 78;
			2767: Pixel = 75;
			2768: Pixel = 74;
			2769: Pixel = 75;
			2770: Pixel = 69;
			2771: Pixel = 73;
			2772: Pixel = 73;
			2773: Pixel = 61;
			2774: Pixel = 127;
			2775: Pixel = 149;
			2776: Pixel = 80;
			2777: Pixel = 68;
			2778: Pixel = 66;
			2779: Pixel = 65;
			2780: Pixel = 68;
			2781: Pixel = 71;
			2782: Pixel = 78;
			2783: Pixel = 81;
			2784: Pixel = 79;
			2785: Pixel = 81;
			2786: Pixel = 78;
			2787: Pixel = 66;
			2788: Pixel = 83;
			2789: Pixel = 78;
			2790: Pixel = 68;
			2791: Pixel = 66;
			2792: Pixel = 83;
			2793: Pixel = 106;
			2794: Pixel = 97;
			2795: Pixel = 99;
			2796: Pixel = 104;
			2797: Pixel = 79;
			2798: Pixel = 50;
			2799: Pixel = 50;
			2800: Pixel = 130;
			2801: Pixel = 126;
			2802: Pixel = 115;
			2803: Pixel = 193;
			2804: Pixel = 206;
			2805: Pixel = 211;
			2806: Pixel = 235;
			2807: Pixel = 226;
			2808: Pixel = 213;
			2809: Pixel = 128;
			2810: Pixel = 128;
			2811: Pixel = 146;
			2812: Pixel = 93;
			2813: Pixel = 83;
			2814: Pixel = 85;
			2815: Pixel = 81;
			2816: Pixel = 77;
			2817: Pixel = 73;
			2818: Pixel = 84;
			2819: Pixel = 110;
			2820: Pixel = 93;
			2821: Pixel = 67;
			2822: Pixel = 54;
			2823: Pixel = 84;
			2824: Pixel = 141;
			2825: Pixel = 70;
			2826: Pixel = 48;
			2827: Pixel = 61;
			2828: Pixel = 71;
			2829: Pixel = 63;
			2830: Pixel = 60;
			2831: Pixel = 77;
			2832: Pixel = 111;
			2833: Pixel = 146;
			2834: Pixel = 187;
			2835: Pixel = 221;
			2836: Pixel = 244;
			2837: Pixel = 236;
			2838: Pixel = 215;
			2839: Pixel = 171;
			2840: Pixel = 168;
			2841: Pixel = 189;
			2842: Pixel = 141;
			2843: Pixel = 188;
			2844: Pixel = 237;
			2845: Pixel = 253;
			2846: Pixel = 235;
			2847: Pixel = 228;
			2848: Pixel = 227;
			2849: Pixel = 237;
			2850: Pixel = 237;
			2851: Pixel = 247;
			2852: Pixel = 245;
			2853: Pixel = 208;
			2854: Pixel = 205;
			2855: Pixel = 245;
			2856: Pixel = 201;
			2857: Pixel = 152;
			2858: Pixel = 146;
			2859: Pixel = 141;
			2860: Pixel = 136;
			2861: Pixel = 98;
			2862: Pixel = 80;
			2863: Pixel = 82;
			2864: Pixel = 79;
			2865: Pixel = 77;
			2866: Pixel = 78;
			2867: Pixel = 76;
			2868: Pixel = 74;
			2869: Pixel = 75;
			2870: Pixel = 68;
			2871: Pixel = 65;
			2872: Pixel = 65;
			2873: Pixel = 62;
			2874: Pixel = 107;
			2875: Pixel = 146;
			2876: Pixel = 80;
			2877: Pixel = 66;
			2878: Pixel = 65;
			2879: Pixel = 68;
			2880: Pixel = 68;
			2881: Pixel = 74;
			2882: Pixel = 80;
			2883: Pixel = 82;
			2884: Pixel = 82;
			2885: Pixel = 84;
			2886: Pixel = 75;
			2887: Pixel = 69;
			2888: Pixel = 84;
			2889: Pixel = 82;
			2890: Pixel = 73;
			2891: Pixel = 67;
			2892: Pixel = 74;
			2893: Pixel = 103;
			2894: Pixel = 100;
			2895: Pixel = 97;
			2896: Pixel = 101;
			2897: Pixel = 84;
			2898: Pixel = 78;
			2899: Pixel = 142;
			2900: Pixel = 78;
			2901: Pixel = 70;
			2902: Pixel = 76;
			2903: Pixel = 189;
			2904: Pixel = 217;
			2905: Pixel = 185;
			2906: Pixel = 222;
			2907: Pixel = 220;
			2908: Pixel = 221;
			2909: Pixel = 143;
			2910: Pixel = 153;
			2911: Pixel = 142;
			2912: Pixel = 102;
			2913: Pixel = 80;
			2914: Pixel = 83;
			2915: Pixel = 80;
			2916: Pixel = 76;
			2917: Pixel = 75;
			2918: Pixel = 77;
			2919: Pixel = 109;
			2920: Pixel = 97;
			2921: Pixel = 75;
			2922: Pixel = 53;
			2923: Pixel = 60;
			2924: Pixel = 65;
			2925: Pixel = 54;
			2926: Pixel = 49;
			2927: Pixel = 55;
			2928: Pixel = 68;
			2929: Pixel = 60;
			2930: Pixel = 53;
			2931: Pixel = 70;
			2932: Pixel = 104;
			2933: Pixel = 144;
			2934: Pixel = 177;
			2935: Pixel = 210;
			2936: Pixel = 241;
			2937: Pixel = 244;
			2938: Pixel = 227;
			2939: Pixel = 161;
			2940: Pixel = 127;
			2941: Pixel = 140;
			2942: Pixel = 186;
			2943: Pixel = 250;
			2944: Pixel = 248;
			2945: Pixel = 246;
			2946: Pixel = 242;
			2947: Pixel = 239;
			2948: Pixel = 233;
			2949: Pixel = 196;
			2950: Pixel = 219;
			2951: Pixel = 251;
			2952: Pixel = 246;
			2953: Pixel = 234;
			2954: Pixel = 223;
			2955: Pixel = 211;
			2956: Pixel = 175;
			2957: Pixel = 151;
			2958: Pixel = 137;
			2959: Pixel = 139;
			2960: Pixel = 126;
			2961: Pixel = 86;
			2962: Pixel = 83;
			2963: Pixel = 81;
			2964: Pixel = 79;
			2965: Pixel = 77;
			2966: Pixel = 76;
			2967: Pixel = 75;
			2968: Pixel = 74;
			2969: Pixel = 75;
			2970: Pixel = 70;
			2971: Pixel = 68;
			2972: Pixel = 89;
			2973: Pixel = 61;
			2974: Pixel = 84;
			2975: Pixel = 117;
			2976: Pixel = 81;
			2977: Pixel = 64;
			2978: Pixel = 63;
			2979: Pixel = 63;
			2980: Pixel = 67;
			2981: Pixel = 74;
			2982: Pixel = 80;
			2983: Pixel = 83;
			2984: Pixel = 84;
			2985: Pixel = 83;
			2986: Pixel = 74;
			2987: Pixel = 75;
			2988: Pixel = 87;
			2989: Pixel = 80;
			2990: Pixel = 75;
			2991: Pixel = 68;
			2992: Pixel = 73;
			2993: Pixel = 93;
			2994: Pixel = 96;
			2995: Pixel = 104;
			2996: Pixel = 131;
			2997: Pixel = 176;
			2998: Pixel = 228;
			2999: Pixel = 255;
			3000: Pixel = 76;
			3001: Pixel = 76;
			3002: Pixel = 76;
			3003: Pixel = 117;
			3004: Pixel = 117;
			3005: Pixel = 83;
			3006: Pixel = 191;
			3007: Pixel = 216;
			3008: Pixel = 218;
			3009: Pixel = 161;
			3010: Pixel = 114;
			3011: Pixel = 112;
			3012: Pixel = 114;
			3013: Pixel = 80;
			3014: Pixel = 83;
			3015: Pixel = 80;
			3016: Pixel = 78;
			3017: Pixel = 75;
			3018: Pixel = 72;
			3019: Pixel = 103;
			3020: Pixel = 103;
			3021: Pixel = 84;
			3022: Pixel = 57;
			3023: Pixel = 53;
			3024: Pixel = 57;
			3025: Pixel = 52;
			3026: Pixel = 47;
			3027: Pixel = 52;
			3028: Pixel = 72;
			3029: Pixel = 64;
			3030: Pixel = 54;
			3031: Pixel = 60;
			3032: Pixel = 94;
			3033: Pixel = 138;
			3034: Pixel = 168;
			3035: Pixel = 198;
			3036: Pixel = 232;
			3037: Pixel = 255;
			3038: Pixel = 205;
			3039: Pixel = 173;
			3040: Pixel = 217;
			3041: Pixel = 219;
			3042: Pixel = 249;
			3043: Pixel = 247;
			3044: Pixel = 246;
			3045: Pixel = 246;
			3046: Pixel = 251;
			3047: Pixel = 221;
			3048: Pixel = 168;
			3049: Pixel = 144;
			3050: Pixel = 218;
			3051: Pixel = 251;
			3052: Pixel = 247;
			3053: Pixel = 241;
			3054: Pixel = 212;
			3055: Pixel = 209;
			3056: Pixel = 222;
			3057: Pixel = 212;
			3058: Pixel = 146;
			3059: Pixel = 129;
			3060: Pixel = 116;
			3061: Pixel = 84;
			3062: Pixel = 83;
			3063: Pixel = 80;
			3064: Pixel = 79;
			3065: Pixel = 76;
			3066: Pixel = 76;
			3067: Pixel = 75;
			3068: Pixel = 73;
			3069: Pixel = 72;
			3070: Pixel = 75;
			3071: Pixel = 70;
			3072: Pixel = 92;
			3073: Pixel = 53;
			3074: Pixel = 67;
			3075: Pixel = 95;
			3076: Pixel = 77;
			3077: Pixel = 61;
			3078: Pixel = 62;
			3079: Pixel = 63;
			3080: Pixel = 68;
			3081: Pixel = 72;
			3082: Pixel = 77;
			3083: Pixel = 78;
			3084: Pixel = 83;
			3085: Pixel = 85;
			3086: Pixel = 74;
			3087: Pixel = 78;
			3088: Pixel = 88;
			3089: Pixel = 81;
			3090: Pixel = 78;
			3091: Pixel = 71;
			3092: Pixel = 64;
			3093: Pixel = 101;
			3094: Pixel = 156;
			3095: Pixel = 213;
			3096: Pixel = 244;
			3097: Pixel = 255;
			3098: Pixel = 250;
			3099: Pixel = 214;
			3100: Pixel = 75;
			3101: Pixel = 78;
			3102: Pixel = 76;
			3103: Pixel = 75;
			3104: Pixel = 82;
			3105: Pixel = 75;
			3106: Pixel = 170;
			3107: Pixel = 220;
			3108: Pixel = 217;
			3109: Pixel = 178;
			3110: Pixel = 114;
			3111: Pixel = 124;
			3112: Pixel = 123;
			3113: Pixel = 83;
			3114: Pixel = 83;
			3115: Pixel = 82;
			3116: Pixel = 80;
			3117: Pixel = 76;
			3118: Pixel = 74;
			3119: Pixel = 87;
			3120: Pixel = 120;
			3121: Pixel = 102;
			3122: Pixel = 63;
			3123: Pixel = 48;
			3124: Pixel = 52;
			3125: Pixel = 49;
			3126: Pixel = 46;
			3127: Pixel = 50;
			3128: Pixel = 67;
			3129: Pixel = 70;
			3130: Pixel = 59;
			3131: Pixel = 56;
			3132: Pixel = 82;
			3133: Pixel = 127;
			3134: Pixel = 159;
			3135: Pixel = 194;
			3136: Pixel = 201;
			3137: Pixel = 165;
			3138: Pixel = 172;
			3139: Pixel = 183;
			3140: Pixel = 250;
			3141: Pixel = 243;
			3142: Pixel = 247;
			3143: Pixel = 247;
			3144: Pixel = 246;
			3145: Pixel = 251;
			3146: Pixel = 215;
			3147: Pixel = 155;
			3148: Pixel = 138;
			3149: Pixel = 149;
			3150: Pixel = 203;
			3151: Pixel = 242;
			3152: Pixel = 247;
			3153: Pixel = 203;
			3154: Pixel = 223;
			3155: Pixel = 250;
			3156: Pixel = 249;
			3157: Pixel = 251;
			3158: Pixel = 203;
			3159: Pixel = 131;
			3160: Pixel = 109;
			3161: Pixel = 86;
			3162: Pixel = 85;
			3163: Pixel = 82;
			3164: Pixel = 79;
			3165: Pixel = 77;
			3166: Pixel = 77;
			3167: Pixel = 75;
			3168: Pixel = 73;
			3169: Pixel = 76;
			3170: Pixel = 75;
			3171: Pixel = 59;
			3172: Pixel = 47;
			3173: Pixel = 49;
			3174: Pixel = 66;
			3175: Pixel = 88;
			3176: Pixel = 72;
			3177: Pixel = 57;
			3178: Pixel = 61;
			3179: Pixel = 66;
			3180: Pixel = 69;
			3181: Pixel = 73;
			3182: Pixel = 75;
			3183: Pixel = 76;
			3184: Pixel = 78;
			3185: Pixel = 80;
			3186: Pixel = 79;
			3187: Pixel = 80;
			3188: Pixel = 78;
			3189: Pixel = 79;
			3190: Pixel = 70;
			3191: Pixel = 75;
			3192: Pixel = 147;
			3193: Pixel = 228;
			3194: Pixel = 244;
			3195: Pixel = 254;
			3196: Pixel = 246;
			3197: Pixel = 210;
			3198: Pixel = 159;
			3199: Pixel = 137;
			3200: Pixel = 74;
			3201: Pixel = 71;
			3202: Pixel = 71;
			3203: Pixel = 73;
			3204: Pixel = 85;
			3205: Pixel = 67;
			3206: Pixel = 141;
			3207: Pixel = 221;
			3208: Pixel = 216;
			3209: Pixel = 195;
			3210: Pixel = 131;
			3211: Pixel = 129;
			3212: Pixel = 127;
			3213: Pixel = 89;
			3214: Pixel = 85;
			3215: Pixel = 82;
			3216: Pixel = 79;
			3217: Pixel = 77;
			3218: Pixel = 76;
			3219: Pixel = 75;
			3220: Pixel = 107;
			3221: Pixel = 101;
			3222: Pixel = 75;
			3223: Pixel = 51;
			3224: Pixel = 47;
			3225: Pixel = 49;
			3226: Pixel = 46;
			3227: Pixel = 48;
			3228: Pixel = 55;
			3229: Pixel = 71;
			3230: Pixel = 67;
			3231: Pixel = 53;
			3232: Pixel = 70;
			3233: Pixel = 115;
			3234: Pixel = 150;
			3235: Pixel = 179;
			3236: Pixel = 211;
			3237: Pixel = 131;
			3238: Pixel = 162;
			3239: Pixel = 237;
			3240: Pixel = 247;
			3241: Pixel = 246;
			3242: Pixel = 246;
			3243: Pixel = 246;
			3244: Pixel = 250;
			3245: Pixel = 215;
			3246: Pixel = 166;
			3247: Pixel = 147;
			3248: Pixel = 133;
			3249: Pixel = 129;
			3250: Pixel = 184;
			3251: Pixel = 225;
			3252: Pixel = 193;
			3253: Pixel = 209;
			3254: Pixel = 255;
			3255: Pixel = 245;
			3256: Pixel = 244;
			3257: Pixel = 225;
			3258: Pixel = 196;
			3259: Pixel = 148;
			3260: Pixel = 112;
			3261: Pixel = 91;
			3262: Pixel = 86;
			3263: Pixel = 83;
			3264: Pixel = 82;
			3265: Pixel = 78;
			3266: Pixel = 75;
			3267: Pixel = 76;
			3268: Pixel = 76;
			3269: Pixel = 77;
			3270: Pixel = 69;
			3271: Pixel = 55;
			3272: Pixel = 51;
			3273: Pixel = 51;
			3274: Pixel = 61;
			3275: Pixel = 81;
			3276: Pixel = 67;
			3277: Pixel = 53;
			3278: Pixel = 58;
			3279: Pixel = 63;
			3280: Pixel = 68;
			3281: Pixel = 72;
			3282: Pixel = 75;
			3283: Pixel = 75;
			3284: Pixel = 73;
			3285: Pixel = 73;
			3286: Pixel = 76;
			3287: Pixel = 97;
			3288: Pixel = 103;
			3289: Pixel = 84;
			3290: Pixel = 135;
			3291: Pixel = 203;
			3292: Pixel = 253;
			3293: Pixel = 255;
			3294: Pixel = 241;
			3295: Pixel = 203;
			3296: Pixel = 176;
			3297: Pixel = 124;
			3298: Pixel = 157;
			3299: Pixel = 202;
			3300: Pixel = 69;
			3301: Pixel = 70;
			3302: Pixel = 72;
			3303: Pixel = 72;
			3304: Pixel = 75;
			3305: Pixel = 69;
			3306: Pixel = 117;
			3307: Pixel = 221;
			3308: Pixel = 216;
			3309: Pixel = 214;
			3310: Pixel = 136;
			3311: Pixel = 120;
			3312: Pixel = 130;
			3313: Pixel = 98;
			3314: Pixel = 82;
			3315: Pixel = 84;
			3316: Pixel = 80;
			3317: Pixel = 76;
			3318: Pixel = 77;
			3319: Pixel = 72;
			3320: Pixel = 85;
			3321: Pixel = 105;
			3322: Pixel = 83;
			3323: Pixel = 62;
			3324: Pixel = 49;
			3325: Pixel = 49;
			3326: Pixel = 48;
			3327: Pixel = 50;
			3328: Pixel = 51;
			3329: Pixel = 62;
			3330: Pixel = 73;
			3331: Pixel = 56;
			3332: Pixel = 56;
			3333: Pixel = 100;
			3334: Pixel = 140;
			3335: Pixel = 166;
			3336: Pixel = 208;
			3337: Pixel = 238;
			3338: Pixel = 238;
			3339: Pixel = 251;
			3340: Pixel = 246;
			3341: Pixel = 247;
			3342: Pixel = 244;
			3343: Pixel = 250;
			3344: Pixel = 226;
			3345: Pixel = 175;
			3346: Pixel = 158;
			3347: Pixel = 131;
			3348: Pixel = 113;
			3349: Pixel = 124;
			3350: Pixel = 162;
			3351: Pixel = 185;
			3352: Pixel = 156;
			3353: Pixel = 237;
			3354: Pixel = 248;
			3355: Pixel = 247;
			3356: Pixel = 240;
			3357: Pixel = 230;
			3358: Pixel = 211;
			3359: Pixel = 162;
			3360: Pixel = 117;
			3361: Pixel = 91;
			3362: Pixel = 87;
			3363: Pixel = 85;
			3364: Pixel = 83;
			3365: Pixel = 79;
			3366: Pixel = 77;
			3367: Pixel = 76;
			3368: Pixel = 76;
			3369: Pixel = 77;
			3370: Pixel = 64;
			3371: Pixel = 49;
			3372: Pixel = 50;
			3373: Pixel = 49;
			3374: Pixel = 60;
			3375: Pixel = 79;
			3376: Pixel = 66;
			3377: Pixel = 54;
			3378: Pixel = 58;
			3379: Pixel = 63;
			3380: Pixel = 67;
			3381: Pixel = 69;
			3382: Pixel = 74;
			3383: Pixel = 75;
			3384: Pixel = 78;
			3385: Pixel = 76;
			3386: Pixel = 73;
			3387: Pixel = 108;
			3388: Pixel = 209;
			3389: Pixel = 212;
			3390: Pixel = 254;
			3391: Pixel = 255;
			3392: Pixel = 233;
			3393: Pixel = 207;
			3394: Pixel = 179;
			3395: Pixel = 135;
			3396: Pixel = 109;
			3397: Pixel = 96;
			3398: Pixel = 198;
			3399: Pixel = 253;
			3400: Pixel = 72;
			3401: Pixel = 75;
			3402: Pixel = 77;
			3403: Pixel = 78;
			3404: Pixel = 79;
			3405: Pixel = 70;
			3406: Pixel = 96;
			3407: Pixel = 224;
			3408: Pixel = 225;
			3409: Pixel = 235;
			3410: Pixel = 153;
			3411: Pixel = 113;
			3412: Pixel = 130;
			3413: Pixel = 104;
			3414: Pixel = 83;
			3415: Pixel = 86;
			3416: Pixel = 83;
			3417: Pixel = 80;
			3418: Pixel = 77;
			3419: Pixel = 76;
			3420: Pixel = 73;
			3421: Pixel = 96;
			3422: Pixel = 91;
			3423: Pixel = 73;
			3424: Pixel = 54;
			3425: Pixel = 49;
			3426: Pixel = 49;
			3427: Pixel = 50;
			3428: Pixel = 52;
			3429: Pixel = 53;
			3430: Pixel = 56;
			3431: Pixel = 57;
			3432: Pixel = 48;
			3433: Pixel = 83;
			3434: Pixel = 128;
			3435: Pixel = 157;
			3436: Pixel = 199;
			3437: Pixel = 239;
			3438: Pixel = 248;
			3439: Pixel = 244;
			3440: Pixel = 247;
			3441: Pixel = 246;
			3442: Pixel = 251;
			3443: Pixel = 232;
			3444: Pixel = 180;
			3445: Pixel = 178;
			3446: Pixel = 168;
			3447: Pixel = 118;
			3448: Pixel = 93;
			3449: Pixel = 170;
			3450: Pixel = 164;
			3451: Pixel = 140;
			3452: Pixel = 149;
			3453: Pixel = 229;
			3454: Pixel = 246;
			3455: Pixel = 250;
			3456: Pixel = 233;
			3457: Pixel = 234;
			3458: Pixel = 245;
			3459: Pixel = 208;
			3460: Pixel = 136;
			3461: Pixel = 89;
			3462: Pixel = 90;
			3463: Pixel = 86;
			3464: Pixel = 85;
			3465: Pixel = 82;
			3466: Pixel = 78;
			3467: Pixel = 78;
			3468: Pixel = 76;
			3469: Pixel = 78;
			3470: Pixel = 63;
			3471: Pixel = 48;
			3472: Pixel = 48;
			3473: Pixel = 48;
			3474: Pixel = 62;
			3475: Pixel = 73;
			3476: Pixel = 64;
			3477: Pixel = 56;
			3478: Pixel = 58;
			3479: Pixel = 61;
			3480: Pixel = 64;
			3481: Pixel = 68;
			3482: Pixel = 74;
			3483: Pixel = 78;
			3484: Pixel = 76;
			3485: Pixel = 75;
			3486: Pixel = 94;
			3487: Pixel = 122;
			3488: Pixel = 232;
			3489: Pixel = 246;
			3490: Pixel = 232;
			3491: Pixel = 200;
			3492: Pixel = 159;
			3493: Pixel = 134;
			3494: Pixel = 123;
			3495: Pixel = 81;
			3496: Pixel = 98;
			3497: Pixel = 108;
			3498: Pixel = 117;
			3499: Pixel = 189;
			3500: Pixel = 78;
			3501: Pixel = 75;
			3502: Pixel = 71;
			3503: Pixel = 75;
			3504: Pixel = 87;
			3505: Pixel = 105;
			3506: Pixel = 138;
			3507: Pixel = 229;
			3508: Pixel = 241;
			3509: Pixel = 254;
			3510: Pixel = 186;
			3511: Pixel = 109;
			3512: Pixel = 124;
			3513: Pixel = 113;
			3514: Pixel = 87;
			3515: Pixel = 90;
			3516: Pixel = 84;
			3517: Pixel = 81;
			3518: Pixel = 78;
			3519: Pixel = 74;
			3520: Pixel = 74;
			3521: Pixel = 74;
			3522: Pixel = 93;
			3523: Pixel = 82;
			3524: Pixel = 67;
			3525: Pixel = 54;
			3526: Pixel = 51;
			3527: Pixel = 50;
			3528: Pixel = 52;
			3529: Pixel = 50;
			3530: Pixel = 62;
			3531: Pixel = 72;
			3532: Pixel = 43;
			3533: Pixel = 65;
			3534: Pixel = 115;
			3535: Pixel = 148;
			3536: Pixel = 196;
			3537: Pixel = 224;
			3538: Pixel = 242;
			3539: Pixel = 230;
			3540: Pixel = 243;
			3541: Pixel = 250;
			3542: Pixel = 243;
			3543: Pixel = 175;
			3544: Pixel = 172;
			3545: Pixel = 189;
			3546: Pixel = 190;
			3547: Pixel = 126;
			3548: Pixel = 96;
			3549: Pixel = 163;
			3550: Pixel = 171;
			3551: Pixel = 120;
			3552: Pixel = 135;
			3553: Pixel = 187;
			3554: Pixel = 234;
			3555: Pixel = 246;
			3556: Pixel = 248;
			3557: Pixel = 250;
			3558: Pixel = 238;
			3559: Pixel = 219;
			3560: Pixel = 180;
			3561: Pixel = 105;
			3562: Pixel = 88;
			3563: Pixel = 88;
			3564: Pixel = 85;
			3565: Pixel = 82;
			3566: Pixel = 81;
			3567: Pixel = 80;
			3568: Pixel = 77;
			3569: Pixel = 74;
			3570: Pixel = 64;
			3571: Pixel = 46;
			3572: Pixel = 42;
			3573: Pixel = 56;
			3574: Pixel = 79;
			3575: Pixel = 88;
			3576: Pixel = 66;
			3577: Pixel = 56;
			3578: Pixel = 59;
			3579: Pixel = 59;
			3580: Pixel = 64;
			3581: Pixel = 69;
			3582: Pixel = 71;
			3583: Pixel = 69;
			3584: Pixel = 81;
			3585: Pixel = 142;
			3586: Pixel = 211;
			3587: Pixel = 199;
			3588: Pixel = 153;
			3589: Pixel = 189;
			3590: Pixel = 148;
			3591: Pixel = 116;
			3592: Pixel = 85;
			3593: Pixel = 71;
			3594: Pixel = 71;
			3595: Pixel = 68;
			3596: Pixel = 110;
			3597: Pixel = 108;
			3598: Pixel = 82;
			3599: Pixel = 106;
			3600: Pixel = 83;
			3601: Pixel = 100;
			3602: Pixel = 133;
			3603: Pixel = 171;
			3604: Pixel = 200;
			3605: Pixel = 205;
			3606: Pixel = 207;
			3607: Pixel = 236;
			3608: Pixel = 248;
			3609: Pixel = 252;
			3610: Pixel = 218;
			3611: Pixel = 116;
			3612: Pixel = 120;
			3613: Pixel = 121;
			3614: Pixel = 90;
			3615: Pixel = 91;
			3616: Pixel = 86;
			3617: Pixel = 82;
			3618: Pixel = 81;
			3619: Pixel = 75;
			3620: Pixel = 75;
			3621: Pixel = 70;
			3622: Pixel = 78;
			3623: Pixel = 92;
			3624: Pixel = 79;
			3625: Pixel = 61;
			3626: Pixel = 52;
			3627: Pixel = 55;
			3628: Pixel = 53;
			3629: Pixel = 51;
			3630: Pixel = 102;
			3631: Pixel = 89;
			3632: Pixel = 48;
			3633: Pixel = 53;
			3634: Pixel = 95;
			3635: Pixel = 139;
			3636: Pixel = 195;
			3637: Pixel = 215;
			3638: Pixel = 223;
			3639: Pixel = 215;
			3640: Pixel = 232;
			3641: Pixel = 247;
			3642: Pixel = 191;
			3643: Pixel = 163;
			3644: Pixel = 170;
			3645: Pixel = 152;
			3646: Pixel = 153;
			3647: Pixel = 111;
			3648: Pixel = 106;
			3649: Pixel = 148;
			3650: Pixel = 140;
			3651: Pixel = 112;
			3652: Pixel = 136;
			3653: Pixel = 207;
			3654: Pixel = 242;
			3655: Pixel = 242;
			3656: Pixel = 247;
			3657: Pixel = 240;
			3658: Pixel = 222;
			3659: Pixel = 231;
			3660: Pixel = 211;
			3661: Pixel = 150;
			3662: Pixel = 91;
			3663: Pixel = 88;
			3664: Pixel = 86;
			3665: Pixel = 85;
			3666: Pixel = 82;
			3667: Pixel = 82;
			3668: Pixel = 79;
			3669: Pixel = 76;
			3670: Pixel = 65;
			3671: Pixel = 50;
			3672: Pixel = 45;
			3673: Pixel = 59;
			3674: Pixel = 95;
			3675: Pixel = 104;
			3676: Pixel = 69;
			3677: Pixel = 59;
			3678: Pixel = 62;
			3679: Pixel = 65;
			3680: Pixel = 62;
			3681: Pixel = 59;
			3682: Pixel = 82;
			3683: Pixel = 146;
			3684: Pixel = 221;
			3685: Pixel = 255;
			3686: Pixel = 206;
			3687: Pixel = 106;
			3688: Pixel = 86;
			3689: Pixel = 124;
			3690: Pixel = 115;
			3691: Pixel = 91;
			3692: Pixel = 76;
			3693: Pixel = 67;
			3694: Pixel = 76;
			3695: Pixel = 78;
			3696: Pixel = 85;
			3697: Pixel = 88;
			3698: Pixel = 63;
			3699: Pixel = 76;
			3700: Pixel = 188;
			3701: Pixel = 223;
			3702: Pixel = 244;
			3703: Pixel = 248;
			3704: Pixel = 237;
			3705: Pixel = 227;
			3706: Pixel = 223;
			3707: Pixel = 238;
			3708: Pixel = 248;
			3709: Pixel = 248;
			3710: Pixel = 241;
			3711: Pixel = 135;
			3712: Pixel = 117;
			3713: Pixel = 125;
			3714: Pixel = 91;
			3715: Pixel = 89;
			3716: Pixel = 86;
			3717: Pixel = 82;
			3718: Pixel = 80;
			3719: Pixel = 78;
			3720: Pixel = 71;
			3721: Pixel = 72;
			3722: Pixel = 68;
			3723: Pixel = 80;
			3724: Pixel = 89;
			3725: Pixel = 75;
			3726: Pixel = 59;
			3727: Pixel = 51;
			3728: Pixel = 54;
			3729: Pixel = 57;
			3730: Pixel = 73;
			3731: Pixel = 91;
			3732: Pixel = 66;
			3733: Pixel = 49;
			3734: Pixel = 76;
			3735: Pixel = 134;
			3736: Pixel = 191;
			3737: Pixel = 207;
			3738: Pixel = 205;
			3739: Pixel = 212;
			3740: Pixel = 224;
			3741: Pixel = 205;
			3742: Pixel = 167;
			3743: Pixel = 154;
			3744: Pixel = 121;
			3745: Pixel = 152;
			3746: Pixel = 185;
			3747: Pixel = 169;
			3748: Pixel = 142;
			3749: Pixel = 153;
			3750: Pixel = 170;
			3751: Pixel = 164;
			3752: Pixel = 219;
			3753: Pixel = 247;
			3754: Pixel = 246;
			3755: Pixel = 244;
			3756: Pixel = 246;
			3757: Pixel = 245;
			3758: Pixel = 245;
			3759: Pixel = 240;
			3760: Pixel = 230;
			3761: Pixel = 197;
			3762: Pixel = 128;
			3763: Pixel = 84;
			3764: Pixel = 88;
			3765: Pixel = 85;
			3766: Pixel = 82;
			3767: Pixel = 83;
			3768: Pixel = 80;
			3769: Pixel = 77;
			3770: Pixel = 66;
			3771: Pixel = 53;
			3772: Pixel = 55;
			3773: Pixel = 81;
			3774: Pixel = 80;
			3775: Pixel = 104;
			3776: Pixel = 92;
			3777: Pixel = 66;
			3778: Pixel = 58;
			3779: Pixel = 58;
			3780: Pixel = 85;
			3781: Pixel = 156;
			3782: Pixel = 230;
			3783: Pixel = 255;
			3784: Pixel = 221;
			3785: Pixel = 159;
			3786: Pixel = 114;
			3787: Pixel = 118;
			3788: Pixel = 118;
			3789: Pixel = 110;
			3790: Pixel = 117;
			3791: Pixel = 116;
			3792: Pixel = 108;
			3793: Pixel = 87;
			3794: Pixel = 78;
			3795: Pixel = 75;
			3796: Pixel = 76;
			3797: Pixel = 81;
			3798: Pixel = 55;
			3799: Pixel = 57;
			3800: Pixel = 219;
			3801: Pixel = 239;
			3802: Pixel = 241;
			3803: Pixel = 238;
			3804: Pixel = 235;
			3805: Pixel = 216;
			3806: Pixel = 213;
			3807: Pixel = 235;
			3808: Pixel = 248;
			3809: Pixel = 246;
			3810: Pixel = 251;
			3811: Pixel = 161;
			3812: Pixel = 115;
			3813: Pixel = 127;
			3814: Pixel = 98;
			3815: Pixel = 87;
			3816: Pixel = 83;
			3817: Pixel = 80;
			3818: Pixel = 79;
			3819: Pixel = 76;
			3820: Pixel = 73;
			3821: Pixel = 71;
			3822: Pixel = 70;
			3823: Pixel = 66;
			3824: Pixel = 75;
			3825: Pixel = 84;
			3826: Pixel = 78;
			3827: Pixel = 67;
			3828: Pixel = 52;
			3829: Pixel = 53;
			3830: Pixel = 56;
			3831: Pixel = 97;
			3832: Pixel = 76;
			3833: Pixel = 52;
			3834: Pixel = 59;
			3835: Pixel = 127;
			3836: Pixel = 193;
			3837: Pixel = 200;
			3838: Pixel = 203;
			3839: Pixel = 208;
			3840: Pixel = 211;
			3841: Pixel = 179;
			3842: Pixel = 162;
			3843: Pixel = 124;
			3844: Pixel = 169;
			3845: Pixel = 223;
			3846: Pixel = 188;
			3847: Pixel = 142;
			3848: Pixel = 157;
			3849: Pixel = 206;
			3850: Pixel = 247;
			3851: Pixel = 214;
			3852: Pixel = 240;
			3853: Pixel = 243;
			3854: Pixel = 245;
			3855: Pixel = 245;
			3856: Pixel = 246;
			3857: Pixel = 247;
			3858: Pixel = 247;
			3859: Pixel = 243;
			3860: Pixel = 232;
			3861: Pixel = 221;
			3862: Pixel = 190;
			3863: Pixel = 116;
			3864: Pixel = 81;
			3865: Pixel = 85;
			3866: Pixel = 84;
			3867: Pixel = 81;
			3868: Pixel = 78;
			3869: Pixel = 76;
			3870: Pixel = 66;
			3871: Pixel = 54;
			3872: Pixel = 56;
			3873: Pixel = 91;
			3874: Pixel = 146;
			3875: Pixel = 156;
			3876: Pixel = 101;
			3877: Pixel = 57;
			3878: Pixel = 92;
			3879: Pixel = 165;
			3880: Pixel = 234;
			3881: Pixel = 255;
			3882: Pixel = 212;
			3883: Pixel = 139;
			3884: Pixel = 88;
			3885: Pixel = 81;
			3886: Pixel = 100;
			3887: Pixel = 128;
			3888: Pixel = 155;
			3889: Pixel = 143;
			3890: Pixel = 117;
			3891: Pixel = 117;
			3892: Pixel = 130;
			3893: Pixel = 117;
			3894: Pixel = 94;
			3895: Pixel = 79;
			3896: Pixel = 76;
			3897: Pixel = 68;
			3898: Pixel = 50;
			3899: Pixel = 47;
			3900: Pixel = 174;
			3901: Pixel = 222;
			3902: Pixel = 236;
			3903: Pixel = 241;
			3904: Pixel = 240;
			3905: Pixel = 217;
			3906: Pixel = 211;
			3907: Pixel = 225;
			3908: Pixel = 248;
			3909: Pixel = 245;
			3910: Pixel = 255;
			3911: Pixel = 185;
			3912: Pixel = 115;
			3913: Pixel = 129;
			3914: Pixel = 105;
			3915: Pixel = 82;
			3916: Pixel = 82;
			3917: Pixel = 78;
			3918: Pixel = 77;
			3919: Pixel = 76;
			3920: Pixel = 73;
			3921: Pixel = 71;
			3922: Pixel = 70;
			3923: Pixel = 69;
			3924: Pixel = 66;
			3925: Pixel = 69;
			3926: Pixel = 82;
			3927: Pixel = 93;
			3928: Pixel = 68;
			3929: Pixel = 56;
			3930: Pixel = 49;
			3931: Pixel = 80;
			3932: Pixel = 85;
			3933: Pixel = 55;
			3934: Pixel = 55;
			3935: Pixel = 121;
			3936: Pixel = 198;
			3937: Pixel = 190;
			3938: Pixel = 197;
			3939: Pixel = 205;
			3940: Pixel = 187;
			3941: Pixel = 170;
			3942: Pixel = 110;
			3943: Pixel = 151;
			3944: Pixel = 207;
			3945: Pixel = 163;
			3946: Pixel = 117;
			3947: Pixel = 152;
			3948: Pixel = 200;
			3949: Pixel = 204;
			3950: Pixel = 173;
			3951: Pixel = 157;
			3952: Pixel = 204;
			3953: Pixel = 243;
			3954: Pixel = 245;
			3955: Pixel = 247;
			3956: Pixel = 246;
			3957: Pixel = 246;
			3958: Pixel = 244;
			3959: Pixel = 237;
			3960: Pixel = 235;
			3961: Pixel = 239;
			3962: Pixel = 219;
			3963: Pixel = 187;
			3964: Pixel = 109;
			3965: Pixel = 77;
			3966: Pixel = 80;
			3967: Pixel = 77;
			3968: Pixel = 77;
			3969: Pixel = 75;
			3970: Pixel = 66;
			3971: Pixel = 57;
			3972: Pixel = 56;
			3973: Pixel = 45;
			3974: Pixel = 84;
			3975: Pixel = 78;
			3976: Pixel = 109;
			3977: Pixel = 175;
			3978: Pixel = 242;
			3979: Pixel = 249;
			3980: Pixel = 197;
			3981: Pixel = 126;
			3982: Pixel = 74;
			3983: Pixel = 57;
			3984: Pixel = 67;
			3985: Pixel = 67;
			3986: Pixel = 72;
			3987: Pixel = 103;
			3988: Pixel = 142;
			3989: Pixel = 156;
			3990: Pixel = 138;
			3991: Pixel = 122;
			3992: Pixel = 130;
			3993: Pixel = 133;
			3994: Pixel = 120;
			3995: Pixel = 98;
			3996: Pixel = 77;
			3997: Pixel = 55;
			3998: Pixel = 53;
			3999: Pixel = 45;
			4000: Pixel = 170;
			4001: Pixel = 197;
			4002: Pixel = 215;
			4003: Pixel = 223;
			4004: Pixel = 213;
			4005: Pixel = 187;
			4006: Pixel = 138;
			4007: Pixel = 149;
			4008: Pixel = 248;
			4009: Pixel = 245;
			4010: Pixel = 253;
			4011: Pixel = 210;
			4012: Pixel = 114;
			4013: Pixel = 123;
			4014: Pixel = 112;
			4015: Pixel = 80;
			4016: Pixel = 79;
			4017: Pixel = 75;
			4018: Pixel = 75;
			4019: Pixel = 76;
			4020: Pixel = 72;
			4021: Pixel = 71;
			4022: Pixel = 71;
			4023: Pixel = 69;
			4024: Pixel = 69;
			4025: Pixel = 66;
			4026: Pixel = 65;
			4027: Pixel = 71;
			4028: Pixel = 81;
			4029: Pixel = 78;
			4030: Pixel = 68;
			4031: Pixel = 62;
			4032: Pixel = 59;
			4033: Pixel = 61;
			4034: Pixel = 53;
			4035: Pixel = 141;
			4036: Pixel = 187;
			4037: Pixel = 173;
			4038: Pixel = 192;
			4039: Pixel = 192;
			4040: Pixel = 172;
			4041: Pixel = 140;
			4042: Pixel = 125;
			4043: Pixel = 181;
			4044: Pixel = 142;
			4045: Pixel = 117;
			4046: Pixel = 162;
			4047: Pixel = 232;
			4048: Pixel = 228;
			4049: Pixel = 186;
			4050: Pixel = 138;
			4051: Pixel = 174;
			4052: Pixel = 214;
			4053: Pixel = 235;
			4054: Pixel = 241;
			4055: Pixel = 248;
			4056: Pixel = 248;
			4057: Pixel = 245;
			4058: Pixel = 245;
			4059: Pixel = 240;
			4060: Pixel = 233;
			4061: Pixel = 203;
			4062: Pixel = 180;
			4063: Pixel = 179;
			4064: Pixel = 164;
			4065: Pixel = 86;
			4066: Pixel = 75;
			4067: Pixel = 75;
			4068: Pixel = 74;
			4069: Pixel = 75;
			4070: Pixel = 67;
			4071: Pixel = 56;
			4072: Pixel = 48;
			4073: Pixel = 52;
			4074: Pixel = 104;
			4075: Pixel = 188;
			4076: Pixel = 244;
			4077: Pixel = 240;
			4078: Pixel = 180;
			4079: Pixel = 116;
			4080: Pixel = 74;
			4081: Pixel = 64;
			4082: Pixel = 63;
			4083: Pixel = 60;
			4084: Pixel = 60;
			4085: Pixel = 58;
			4086: Pixel = 57;
			4087: Pixel = 76;
			4088: Pixel = 115;
			4089: Pixel = 145;
			4090: Pixel = 153;
			4091: Pixel = 143;
			4092: Pixel = 130;
			4093: Pixel = 133;
			4094: Pixel = 119;
			4095: Pixel = 86;
			4096: Pixel = 55;
			4097: Pixel = 51;
			4098: Pixel = 50;
			4099: Pixel = 45;
			4100: Pixel = 190;
			4101: Pixel = 195;
			4102: Pixel = 203;
			4103: Pixel = 212;
			4104: Pixel = 203;
			4105: Pixel = 115;
			4106: Pixel = 106;
			4107: Pixel = 118;
			4108: Pixel = 227;
			4109: Pixel = 250;
			4110: Pixel = 249;
			4111: Pixel = 226;
			4112: Pixel = 120;
			4113: Pixel = 117;
			4114: Pixel = 119;
			4115: Pixel = 84;
			4116: Pixel = 79;
			4117: Pixel = 76;
			4118: Pixel = 76;
			4119: Pixel = 75;
			4120: Pixel = 72;
			4121: Pixel = 72;
			4122: Pixel = 71;
			4123: Pixel = 71;
			4124: Pixel = 71;
			4125: Pixel = 69;
			4126: Pixel = 67;
			4127: Pixel = 63;
			4128: Pixel = 63;
			4129: Pixel = 68;
			4130: Pixel = 73;
			4131: Pixel = 70;
			4132: Pixel = 68;
			4133: Pixel = 64;
			4134: Pixel = 73;
			4135: Pixel = 200;
			4136: Pixel = 177;
			4137: Pixel = 175;
			4138: Pixel = 184;
			4139: Pixel = 172;
			4140: Pixel = 153;
			4141: Pixel = 116;
			4142: Pixel = 161;
			4143: Pixel = 137;
			4144: Pixel = 135;
			4145: Pixel = 195;
			4146: Pixel = 247;
			4147: Pixel = 240;
			4148: Pixel = 214;
			4149: Pixel = 226;
			4150: Pixel = 212;
			4151: Pixel = 233;
			4152: Pixel = 246;
			4153: Pixel = 227;
			4154: Pixel = 236;
			4155: Pixel = 241;
			4156: Pixel = 241;
			4157: Pixel = 243;
			4158: Pixel = 241;
			4159: Pixel = 216;
			4160: Pixel = 199;
			4161: Pixel = 185;
			4162: Pixel = 174;
			4163: Pixel = 159;
			4164: Pixel = 184;
			4165: Pixel = 118;
			4166: Pixel = 75;
			4167: Pixel = 80;
			4168: Pixel = 79;
			4169: Pixel = 71;
			4170: Pixel = 55;
			4171: Pixel = 63;
			4172: Pixel = 126;
			4173: Pixel = 203;
			4174: Pixel = 250;
			4175: Pixel = 231;
			4176: Pixel = 165;
			4177: Pixel = 99;
			4178: Pixel = 69;
			4179: Pixel = 70;
			4180: Pixel = 73;
			4181: Pixel = 72;
			4182: Pixel = 61;
			4183: Pixel = 53;
			4184: Pixel = 54;
			4185: Pixel = 54;
			4186: Pixel = 60;
			4187: Pixel = 70;
			4188: Pixel = 89;
			4189: Pixel = 123;
			4190: Pixel = 143;
			4191: Pixel = 150;
			4192: Pixel = 141;
			4193: Pixel = 129;
			4194: Pixel = 121;
			4195: Pixel = 103;
			4196: Pixel = 69;
			4197: Pixel = 52;
			4198: Pixel = 52;
			4199: Pixel = 50;
			4200: Pixel = 203;
			4201: Pixel = 209;
			4202: Pixel = 217;
			4203: Pixel = 227;
			4204: Pixel = 240;
			4205: Pixel = 161;
			4206: Pixel = 105;
			4207: Pixel = 119;
			4208: Pixel = 212;
			4209: Pixel = 253;
			4210: Pixel = 248;
			4211: Pixel = 236;
			4212: Pixel = 129;
			4213: Pixel = 112;
			4214: Pixel = 122;
			4215: Pixel = 89;
			4216: Pixel = 81;
			4217: Pixel = 75;
			4218: Pixel = 74;
			4219: Pixel = 73;
			4220: Pixel = 71;
			4221: Pixel = 71;
			4222: Pixel = 74;
			4223: Pixel = 71;
			4224: Pixel = 70;
			4225: Pixel = 69;
			4226: Pixel = 67;
			4227: Pixel = 67;
			4228: Pixel = 66;
			4229: Pixel = 59;
			4230: Pixel = 54;
			4231: Pixel = 59;
			4232: Pixel = 61;
			4233: Pixel = 52;
			4234: Pixel = 111;
			4235: Pixel = 232;
			4236: Pixel = 166;
			4237: Pixel = 175;
			4238: Pixel = 182;
			4239: Pixel = 154;
			4240: Pixel = 122;
			4241: Pixel = 127;
			4242: Pixel = 137;
			4243: Pixel = 139;
			4244: Pixel = 222;
			4245: Pixel = 249;
			4246: Pixel = 255;
			4247: Pixel = 193;
			4248: Pixel = 122;
			4249: Pixel = 236;
			4250: Pixel = 220;
			4251: Pixel = 218;
			4252: Pixel = 192;
			4253: Pixel = 186;
			4254: Pixel = 218;
			4255: Pixel = 235;
			4256: Pixel = 239;
			4257: Pixel = 228;
			4258: Pixel = 202;
			4259: Pixel = 196;
			4260: Pixel = 186;
			4261: Pixel = 185;
			4262: Pixel = 193;
			4263: Pixel = 159;
			4264: Pixel = 176;
			4265: Pixel = 144;
			4266: Pixel = 84;
			4267: Pixel = 76;
			4268: Pixel = 68;
			4269: Pixel = 86;
			4270: Pixel = 141;
			4271: Pixel = 214;
			4272: Pixel = 254;
			4273: Pixel = 221;
			4274: Pixel = 156;
			4275: Pixel = 96;
			4276: Pixel = 63;
			4277: Pixel = 65;
			4278: Pixel = 70;
			4279: Pixel = 77;
			4280: Pixel = 72;
			4281: Pixel = 68;
			4282: Pixel = 58;
			4283: Pixel = 47;
			4284: Pixel = 46;
			4285: Pixel = 56;
			4286: Pixel = 56;
			4287: Pixel = 60;
			4288: Pixel = 74;
			4289: Pixel = 95;
			4290: Pixel = 118;
			4291: Pixel = 137;
			4292: Pixel = 139;
			4293: Pixel = 127;
			4294: Pixel = 120;
			4295: Pixel = 114;
			4296: Pixel = 90;
			4297: Pixel = 65;
			4298: Pixel = 51;
			4299: Pixel = 51;
			4300: Pixel = 224;
			4301: Pixel = 232;
			4302: Pixel = 240;
			4303: Pixel = 244;
			4304: Pixel = 249;
			4305: Pixel = 235;
			4306: Pixel = 204;
			4307: Pixel = 230;
			4308: Pixel = 244;
			4309: Pixel = 244;
			4310: Pixel = 244;
			4311: Pixel = 237;
			4312: Pixel = 141;
			4313: Pixel = 110;
			4314: Pixel = 119;
			4315: Pixel = 93;
			4316: Pixel = 80;
			4317: Pixel = 77;
			4318: Pixel = 75;
			4319: Pixel = 72;
			4320: Pixel = 70;
			4321: Pixel = 71;
			4322: Pixel = 74;
			4323: Pixel = 73;
			4324: Pixel = 71;
			4325: Pixel = 67;
			4326: Pixel = 66;
			4327: Pixel = 65;
			4328: Pixel = 61;
			4329: Pixel = 58;
			4330: Pixel = 53;
			4331: Pixel = 55;
			4332: Pixel = 57;
			4333: Pixel = 48;
			4334: Pixel = 143;
			4335: Pixel = 229;
			4336: Pixel = 174;
			4337: Pixel = 167;
			4338: Pixel = 170;
			4339: Pixel = 144;
			4340: Pixel = 122;
			4341: Pixel = 130;
			4342: Pixel = 133;
			4343: Pixel = 225;
			4344: Pixel = 252;
			4345: Pixel = 244;
			4346: Pixel = 250;
			4347: Pixel = 230;
			4348: Pixel = 171;
			4349: Pixel = 234;
			4350: Pixel = 220;
			4351: Pixel = 197;
			4352: Pixel = 182;
			4353: Pixel = 183;
			4354: Pixel = 212;
			4355: Pixel = 238;
			4356: Pixel = 206;
			4357: Pixel = 196;
			4358: Pixel = 187;
			4359: Pixel = 186;
			4360: Pixel = 181;
			4361: Pixel = 172;
			4362: Pixel = 140;
			4363: Pixel = 175;
			4364: Pixel = 171;
			4365: Pixel = 134;
			4366: Pixel = 80;
			4367: Pixel = 106;
			4368: Pixel = 164;
			4369: Pixel = 229;
			4370: Pixel = 253;
			4371: Pixel = 213;
			4372: Pixel = 136;
			4373: Pixel = 78;
			4374: Pixel = 73;
			4375: Pixel = 75;
			4376: Pixel = 69;
			4377: Pixel = 70;
			4378: Pixel = 71;
			4379: Pixel = 73;
			4380: Pixel = 74;
			4381: Pixel = 69;
			4382: Pixel = 60;
			4383: Pixel = 45;
			4384: Pixel = 46;
			4385: Pixel = 46;
			4386: Pixel = 50;
			4387: Pixel = 57;
			4388: Pixel = 65;
			4389: Pixel = 74;
			4390: Pixel = 89;
			4391: Pixel = 113;
			4392: Pixel = 126;
			4393: Pixel = 121;
			4394: Pixel = 121;
			4395: Pixel = 113;
			4396: Pixel = 96;
			4397: Pixel = 80;
			4398: Pixel = 57;
			4399: Pixel = 54;
			4400: Pixel = 244;
			4401: Pixel = 247;
			4402: Pixel = 247;
			4403: Pixel = 248;
			4404: Pixel = 247;
			4405: Pixel = 249;
			4406: Pixel = 254;
			4407: Pixel = 250;
			4408: Pixel = 247;
			4409: Pixel = 229;
			4410: Pixel = 230;
			4411: Pixel = 230;
			4412: Pixel = 156;
			4413: Pixel = 110;
			4414: Pixel = 118;
			4415: Pixel = 101;
			4416: Pixel = 80;
			4417: Pixel = 81;
			4418: Pixel = 76;
			4419: Pixel = 75;
			4420: Pixel = 73;
			4421: Pixel = 72;
			4422: Pixel = 71;
			4423: Pixel = 71;
			4424: Pixel = 69;
			4425: Pixel = 67;
			4426: Pixel = 61;
			4427: Pixel = 58;
			4428: Pixel = 57;
			4429: Pixel = 54;
			4430: Pixel = 54;
			4431: Pixel = 56;
			4432: Pixel = 57;
			4433: Pixel = 50;
			4434: Pixel = 126;
			4435: Pixel = 217;
			4436: Pixel = 184;
			4437: Pixel = 160;
			4438: Pixel = 155;
			4439: Pixel = 132;
			4440: Pixel = 126;
			4441: Pixel = 148;
			4442: Pixel = 224;
			4443: Pixel = 252;
			4444: Pixel = 244;
			4445: Pixel = 247;
			4446: Pixel = 246;
			4447: Pixel = 252;
			4448: Pixel = 225;
			4449: Pixel = 209;
			4450: Pixel = 227;
			4451: Pixel = 229;
			4452: Pixel = 234;
			4453: Pixel = 233;
			4454: Pixel = 227;
			4455: Pixel = 184;
			4456: Pixel = 184;
			4457: Pixel = 200;
			4458: Pixel = 184;
			4459: Pixel = 177;
			4460: Pixel = 181;
			4461: Pixel = 174;
			4462: Pixel = 153;
			4463: Pixel = 171;
			4464: Pixel = 170;
			4465: Pixel = 137;
			4466: Pixel = 180;
			4467: Pixel = 244;
			4468: Pixel = 254;
			4469: Pixel = 203;
			4470: Pixel = 131;
			4471: Pixel = 72;
			4472: Pixel = 47;
			4473: Pixel = 54;
			4474: Pixel = 74;
			4475: Pixel = 78;
			4476: Pixel = 67;
			4477: Pixel = 71;
			4478: Pixel = 70;
			4479: Pixel = 73;
			4480: Pixel = 73;
			4481: Pixel = 68;
			4482: Pixel = 64;
			4483: Pixel = 45;
			4484: Pixel = 45;
			4485: Pixel = 43;
			4486: Pixel = 51;
			4487: Pixel = 55;
			4488: Pixel = 62;
			4489: Pixel = 65;
			4490: Pixel = 76;
			4491: Pixel = 91;
			4492: Pixel = 101;
			4493: Pixel = 116;
			4494: Pixel = 121;
			4495: Pixel = 113;
			4496: Pixel = 95;
			4497: Pixel = 79;
			4498: Pixel = 61;
			4499: Pixel = 58;
			4500: Pixel = 247;
			4501: Pixel = 247;
			4502: Pixel = 247;
			4503: Pixel = 247;
			4504: Pixel = 247;
			4505: Pixel = 246;
			4506: Pixel = 245;
			4507: Pixel = 247;
			4508: Pixel = 234;
			4509: Pixel = 211;
			4510: Pixel = 215;
			4511: Pixel = 218;
			4512: Pixel = 162;
			4513: Pixel = 111;
			4514: Pixel = 116;
			4515: Pixel = 107;
			4516: Pixel = 86;
			4517: Pixel = 83;
			4518: Pixel = 75;
			4519: Pixel = 79;
			4520: Pixel = 77;
			4521: Pixel = 70;
			4522: Pixel = 73;
			4523: Pixel = 64;
			4524: Pixel = 59;
			4525: Pixel = 58;
			4526: Pixel = 52;
			4527: Pixel = 54;
			4528: Pixel = 51;
			4529: Pixel = 55;
			4530: Pixel = 59;
			4531: Pixel = 59;
			4532: Pixel = 58;
			4533: Pixel = 51;
			4534: Pixel = 91;
			4535: Pixel = 187;
			4536: Pixel = 150;
			4537: Pixel = 176;
			4538: Pixel = 150;
			4539: Pixel = 119;
			4540: Pixel = 168;
			4541: Pixel = 240;
			4542: Pixel = 252;
			4543: Pixel = 245;
			4544: Pixel = 246;
			4545: Pixel = 247;
			4546: Pixel = 247;
			4547: Pixel = 247;
			4548: Pixel = 242;
			4549: Pixel = 216;
			4550: Pixel = 242;
			4551: Pixel = 246;
			4552: Pixel = 236;
			4553: Pixel = 212;
			4554: Pixel = 185;
			4555: Pixel = 179;
			4556: Pixel = 150;
			4557: Pixel = 165;
			4558: Pixel = 200;
			4559: Pixel = 190;
			4560: Pixel = 168;
			4561: Pixel = 179;
			4562: Pixel = 179;
			4563: Pixel = 168;
			4564: Pixel = 199;
			4565: Pixel = 246;
			4566: Pixel = 249;
			4567: Pixel = 195;
			4568: Pixel = 127;
			4569: Pixel = 82;
			4570: Pixel = 65;
			4571: Pixel = 59;
			4572: Pixel = 55;
			4573: Pixel = 58;
			4574: Pixel = 71;
			4575: Pixel = 73;
			4576: Pixel = 67;
			4577: Pixel = 71;
			4578: Pixel = 68;
			4579: Pixel = 70;
			4580: Pixel = 71;
			4581: Pixel = 67;
			4582: Pixel = 67;
			4583: Pixel = 48;
			4584: Pixel = 44;
			4585: Pixel = 44;
			4586: Pixel = 48;
			4587: Pixel = 53;
			4588: Pixel = 57;
			4589: Pixel = 62;
			4590: Pixel = 66;
			4591: Pixel = 73;
			4592: Pixel = 86;
			4593: Pixel = 102;
			4594: Pixel = 110;
			4595: Pixel = 108;
			4596: Pixel = 91;
			4597: Pixel = 77;
			4598: Pixel = 58;
			4599: Pixel = 67;
			4600: Pixel = 247;
			4601: Pixel = 246;
			4602: Pixel = 247;
			4603: Pixel = 247;
			4604: Pixel = 247;
			4605: Pixel = 247;
			4606: Pixel = 249;
			4607: Pixel = 237;
			4608: Pixel = 206;
			4609: Pixel = 201;
			4610: Pixel = 204;
			4611: Pixel = 207;
			4612: Pixel = 164;
			4613: Pixel = 113;
			4614: Pixel = 116;
			4615: Pixel = 113;
			4616: Pixel = 90;
			4617: Pixel = 83;
			4618: Pixel = 71;
			4619: Pixel = 72;
			4620: Pixel = 73;
			4621: Pixel = 68;
			4622: Pixel = 69;
			4623: Pixel = 65;
			4624: Pixel = 60;
			4625: Pixel = 59;
			4626: Pixel = 56;
			4627: Pixel = 55;
			4628: Pixel = 57;
			4629: Pixel = 67;
			4630: Pixel = 57;
			4631: Pixel = 58;
			4632: Pixel = 60;
			4633: Pixel = 59;
			4634: Pixel = 77;
			4635: Pixel = 136;
			4636: Pixel = 164;
			4637: Pixel = 213;
			4638: Pixel = 139;
			4639: Pixel = 182;
			4640: Pixel = 249;
			4641: Pixel = 249;
			4642: Pixel = 245;
			4643: Pixel = 246;
			4644: Pixel = 247;
			4645: Pixel = 247;
			4646: Pixel = 247;
			4647: Pixel = 247;
			4648: Pixel = 246;
			4649: Pixel = 249;
			4650: Pixel = 250;
			4651: Pixel = 226;
			4652: Pixel = 192;
			4653: Pixel = 188;
			4654: Pixel = 177;
			4655: Pixel = 165;
			4656: Pixel = 113;
			4657: Pixel = 136;
			4658: Pixel = 177;
			4659: Pixel = 171;
			4660: Pixel = 181;
			4661: Pixel = 170;
			4662: Pixel = 163;
			4663: Pixel = 163;
			4664: Pixel = 211;
			4665: Pixel = 193;
			4666: Pixel = 123;
			4667: Pixel = 84;
			4668: Pixel = 76;
			4669: Pixel = 75;
			4670: Pixel = 73;
			4671: Pixel = 61;
			4672: Pixel = 55;
			4673: Pixel = 56;
			4674: Pixel = 71;
			4675: Pixel = 71;
			4676: Pixel = 68;
			4677: Pixel = 70;
			4678: Pixel = 71;
			4679: Pixel = 72;
			4680: Pixel = 68;
			4681: Pixel = 68;
			4682: Pixel = 67;
			4683: Pixel = 57;
			4684: Pixel = 44;
			4685: Pixel = 42;
			4686: Pixel = 48;
			4687: Pixel = 51;
			4688: Pixel = 56;
			4689: Pixel = 58;
			4690: Pixel = 60;
			4691: Pixel = 63;
			4692: Pixel = 74;
			4693: Pixel = 82;
			4694: Pixel = 93;
			4695: Pixel = 97;
			4696: Pixel = 88;
			4697: Pixel = 67;
			4698: Pixel = 72;
			4699: Pixel = 123;
			4700: Pixel = 247;
			4701: Pixel = 247;
			4702: Pixel = 247;
			4703: Pixel = 247;
			4704: Pixel = 247;
			4705: Pixel = 247;
			4706: Pixel = 244;
			4707: Pixel = 218;
			4708: Pixel = 186;
			4709: Pixel = 189;
			4710: Pixel = 201;
			4711: Pixel = 200;
			4712: Pixel = 160;
			4713: Pixel = 119;
			4714: Pixel = 123;
			4715: Pixel = 127;
			4716: Pixel = 92;
			4717: Pixel = 80;
			4718: Pixel = 70;
			4719: Pixel = 67;
			4720: Pixel = 62;
			4721: Pixel = 64;
			4722: Pixel = 64;
			4723: Pixel = 68;
			4724: Pixel = 66;
			4725: Pixel = 65;
			4726: Pixel = 60;
			4727: Pixel = 60;
			4728: Pixel = 65;
			4729: Pixel = 69;
			4730: Pixel = 67;
			4731: Pixel = 75;
			4732: Pixel = 94;
			4733: Pixel = 98;
			4734: Pixel = 93;
			4735: Pixel = 114;
			4736: Pixel = 197;
			4737: Pixel = 210;
			4738: Pixel = 181;
			4739: Pixel = 253;
			4740: Pixel = 247;
			4741: Pixel = 246;
			4742: Pixel = 247;
			4743: Pixel = 247;
			4744: Pixel = 247;
			4745: Pixel = 247;
			4746: Pixel = 247;
			4747: Pixel = 246;
			4748: Pixel = 249;
			4749: Pixel = 245;
			4750: Pixel = 211;
			4751: Pixel = 187;
			4752: Pixel = 185;
			4753: Pixel = 179;
			4754: Pixel = 161;
			4755: Pixel = 146;
			4756: Pixel = 127;
			4757: Pixel = 108;
			4758: Pixel = 116;
			4759: Pixel = 138;
			4760: Pixel = 158;
			4761: Pixel = 165;
			4762: Pixel = 164;
			4763: Pixel = 183;
			4764: Pixel = 172;
			4765: Pixel = 104;
			4766: Pixel = 79;
			4767: Pixel = 85;
			4768: Pixel = 81;
			4769: Pixel = 75;
			4770: Pixel = 68;
			4771: Pixel = 58;
			4772: Pixel = 50;
			4773: Pixel = 54;
			4774: Pixel = 69;
			4775: Pixel = 70;
			4776: Pixel = 66;
			4777: Pixel = 69;
			4778: Pixel = 74;
			4779: Pixel = 71;
			4780: Pixel = 63;
			4781: Pixel = 66;
			4782: Pixel = 72;
			4783: Pixel = 65;
			4784: Pixel = 52;
			4785: Pixel = 44;
			4786: Pixel = 41;
			4787: Pixel = 49;
			4788: Pixel = 51;
			4789: Pixel = 51;
			4790: Pixel = 56;
			4791: Pixel = 59;
			4792: Pixel = 64;
			4793: Pixel = 64;
			4794: Pixel = 72;
			4795: Pixel = 82;
			4796: Pixel = 81;
			4797: Pixel = 55;
			4798: Pixel = 112;
			4799: Pixel = 221;
			4800: Pixel = 247;
			4801: Pixel = 248;
			4802: Pixel = 248;
			4803: Pixel = 247;
			4804: Pixel = 247;
			4805: Pixel = 243;
			4806: Pixel = 228;
			4807: Pixel = 207;
			4808: Pixel = 172;
			4809: Pixel = 169;
			4810: Pixel = 187;
			4811: Pixel = 192;
			4812: Pixel = 155;
			4813: Pixel = 117;
			4814: Pixel = 149;
			4815: Pixel = 137;
			4816: Pixel = 91;
			4817: Pixel = 81;
			4818: Pixel = 80;
			4819: Pixel = 71;
			4820: Pixel = 65;
			4821: Pixel = 63;
			4822: Pixel = 65;
			4823: Pixel = 68;
			4824: Pixel = 68;
			4825: Pixel = 67;
			4826: Pixel = 66;
			4827: Pixel = 81;
			4828: Pixel = 91;
			4829: Pixel = 117;
			4830: Pixel = 135;
			4831: Pixel = 122;
			4832: Pixel = 106;
			4833: Pixel = 91;
			4834: Pixel = 71;
			4835: Pixel = 90;
			4836: Pixel = 194;
			4837: Pixel = 225;
			4838: Pixel = 225;
			4839: Pixel = 244;
			4840: Pixel = 247;
			4841: Pixel = 247;
			4842: Pixel = 247;
			4843: Pixel = 247;
			4844: Pixel = 247;
			4845: Pixel = 247;
			4846: Pixel = 246;
			4847: Pixel = 249;
			4848: Pixel = 240;
			4849: Pixel = 202;
			4850: Pixel = 188;
			4851: Pixel = 189;
			4852: Pixel = 172;
			4853: Pixel = 146;
			4854: Pixel = 153;
			4855: Pixel = 129;
			4856: Pixel = 107;
			4857: Pixel = 110;
			4858: Pixel = 151;
			4859: Pixel = 155;
			4860: Pixel = 136;
			4861: Pixel = 157;
			4862: Pixel = 171;
			4863: Pixel = 186;
			4864: Pixel = 186;
			4865: Pixel = 148;
			4866: Pixel = 87;
			4867: Pixel = 80;
			4868: Pixel = 77;
			4869: Pixel = 75;
			4870: Pixel = 69;
			4871: Pixel = 56;
			4872: Pixel = 49;
			4873: Pixel = 53;
			4874: Pixel = 68;
			4875: Pixel = 67;
			4876: Pixel = 66;
			4877: Pixel = 69;
			4878: Pixel = 72;
			4879: Pixel = 70;
			4880: Pixel = 64;
			4881: Pixel = 66;
			4882: Pixel = 73;
			4883: Pixel = 66;
			4884: Pixel = 56;
			4885: Pixel = 54;
			4886: Pixel = 47;
			4887: Pixel = 45;
			4888: Pixel = 52;
			4889: Pixel = 54;
			4890: Pixel = 54;
			4891: Pixel = 53;
			4892: Pixel = 56;
			4893: Pixel = 60;
			4894: Pixel = 63;
			4895: Pixel = 68;
			4896: Pixel = 60;
			4897: Pixel = 47;
			4898: Pixel = 111;
			4899: Pixel = 228;
			4900: Pixel = 245;
			4901: Pixel = 243;
			4902: Pixel = 242;
			4903: Pixel = 245;
			4904: Pixel = 240;
			4905: Pixel = 231;
			4906: Pixel = 216;
			4907: Pixel = 200;
			4908: Pixel = 163;
			4909: Pixel = 148;
			4910: Pixel = 172;
			4911: Pixel = 180;
			4912: Pixel = 141;
			4913: Pixel = 118;
			4914: Pixel = 117;
			4915: Pixel = 101;
			4916: Pixel = 99;
			4917: Pixel = 86;
			4918: Pixel = 90;
			4919: Pixel = 72;
			4920: Pixel = 68;
			4921: Pixel = 66;
			4922: Pixel = 76;
			4923: Pixel = 81;
			4924: Pixel = 96;
			4925: Pixel = 106;
			4926: Pixel = 125;
			4927: Pixel = 139;
			4928: Pixel = 148;
			4929: Pixel = 141;
			4930: Pixel = 114;
			4931: Pixel = 90;
			4932: Pixel = 76;
			4933: Pixel = 67;
			4934: Pixel = 58;
			4935: Pixel = 64;
			4936: Pixel = 168;
			4937: Pixel = 222;
			4938: Pixel = 162;
			4939: Pixel = 222;
			4940: Pixel = 253;
			4941: Pixel = 246;
			4942: Pixel = 247;
			4943: Pixel = 247;
			4944: Pixel = 247;
			4945: Pixel = 246;
			4946: Pixel = 251;
			4947: Pixel = 231;
			4948: Pixel = 195;
			4949: Pixel = 198;
			4950: Pixel = 182;
			4951: Pixel = 115;
			4952: Pixel = 143;
			4953: Pixel = 145;
			4954: Pixel = 119;
			4955: Pixel = 103;
			4956: Pixel = 108;
			4957: Pixel = 114;
			4958: Pixel = 124;
			4959: Pixel = 142;
			4960: Pixel = 146;
			4961: Pixel = 151;
			4962: Pixel = 165;
			4963: Pixel = 167;
			4964: Pixel = 175;
			4965: Pixel = 176;
			4966: Pixel = 116;
			4967: Pixel = 72;
			4968: Pixel = 75;
			4969: Pixel = 72;
			4970: Pixel = 67;
			4971: Pixel = 57;
			4972: Pixel = 50;
			4973: Pixel = 53;
			4974: Pixel = 67;
			4975: Pixel = 66;
			4976: Pixel = 59;
			4977: Pixel = 64;
			4978: Pixel = 72;
			4979: Pixel = 68;
			4980: Pixel = 64;
			4981: Pixel = 66;
			4982: Pixel = 74;
			4983: Pixel = 69;
			4984: Pixel = 56;
			4985: Pixel = 53;
			4986: Pixel = 56;
			4987: Pixel = 50;
			4988: Pixel = 50;
			4989: Pixel = 53;
			4990: Pixel = 47;
			4991: Pixel = 53;
			4992: Pixel = 54;
			4993: Pixel = 53;
			4994: Pixel = 51;
			4995: Pixel = 68;
			4996: Pixel = 105;
			4997: Pixel = 160;
			4998: Pixel = 217;
			4999: Pixel = 200;
			5000: Pixel = 223;
			5001: Pixel = 222;
			5002: Pixel = 224;
			5003: Pixel = 228;
			5004: Pixel = 222;
			5005: Pixel = 216;
			5006: Pixel = 202;
			5007: Pixel = 179;
			5008: Pixel = 140;
			5009: Pixel = 118;
			5010: Pixel = 151;
			5011: Pixel = 164;
			5012: Pixel = 131;
			5013: Pixel = 111;
			5014: Pixel = 131;
			5015: Pixel = 123;
			5016: Pixel = 121;
			5017: Pixel = 116;
			5018: Pixel = 124;
			5019: Pixel = 107;
			5020: Pixel = 114;
			5021: Pixel = 125;
			5022: Pixel = 139;
			5023: Pixel = 155;
			5024: Pixel = 162;
			5025: Pixel = 164;
			5026: Pixel = 147;
			5027: Pixel = 130;
			5028: Pixel = 115;
			5029: Pixel = 107;
			5030: Pixel = 85;
			5031: Pixel = 69;
			5032: Pixel = 64;
			5033: Pixel = 58;
			5034: Pixel = 57;
			5035: Pixel = 52;
			5036: Pixel = 137;
			5037: Pixel = 186;
			5038: Pixel = 99;
			5039: Pixel = 180;
			5040: Pixel = 255;
			5041: Pixel = 245;
			5042: Pixel = 247;
			5043: Pixel = 246;
			5044: Pixel = 247;
			5045: Pixel = 248;
			5046: Pixel = 218;
			5047: Pixel = 192;
			5048: Pixel = 200;
			5049: Pixel = 184;
			5050: Pixel = 165;
			5051: Pixel = 179;
			5052: Pixel = 119;
			5053: Pixel = 102;
			5054: Pixel = 101;
			5055: Pixel = 96;
			5056: Pixel = 97;
			5057: Pixel = 96;
			5058: Pixel = 107;
			5059: Pixel = 129;
			5060: Pixel = 141;
			5061: Pixel = 146;
			5062: Pixel = 167;
			5063: Pixel = 144;
			5064: Pixel = 157;
			5065: Pixel = 190;
			5066: Pixel = 169;
			5067: Pixel = 94;
			5068: Pixel = 70;
			5069: Pixel = 72;
			5070: Pixel = 66;
			5071: Pixel = 56;
			5072: Pixel = 50;
			5073: Pixel = 53;
			5074: Pixel = 67;
			5075: Pixel = 62;
			5076: Pixel = 84;
			5077: Pixel = 70;
			5078: Pixel = 72;
			5079: Pixel = 70;
			5080: Pixel = 65;
			5081: Pixel = 66;
			5082: Pixel = 68;
			5083: Pixel = 62;
			5084: Pixel = 52;
			5085: Pixel = 58;
			5086: Pixel = 64;
			5087: Pixel = 64;
			5088: Pixel = 59;
			5089: Pixel = 47;
			5090: Pixel = 50;
			5091: Pixel = 46;
			5092: Pixel = 49;
			5093: Pixel = 79;
			5094: Pixel = 140;
			5095: Pixel = 208;
			5096: Pixel = 246;
			5097: Pixel = 230;
			5098: Pixel = 158;
			5099: Pixel = 99;
			5100: Pixel = 205;
			5101: Pixel = 209;
			5102: Pixel = 208;
			5103: Pixel = 206;
			5104: Pixel = 202;
			5105: Pixel = 195;
			5106: Pixel = 174;
			5107: Pixel = 146;
			5108: Pixel = 129;
			5109: Pixel = 146;
			5110: Pixel = 157;
			5111: Pixel = 132;
			5112: Pixel = 125;
			5113: Pixel = 127;
			5114: Pixel = 136;
			5115: Pixel = 134;
			5116: Pixel = 132;
			5117: Pixel = 141;
			5118: Pixel = 146;
			5119: Pixel = 132;
			5120: Pixel = 140;
			5121: Pixel = 146;
			5122: Pixel = 151;
			5123: Pixel = 150;
			5124: Pixel = 128;
			5125: Pixel = 117;
			5126: Pixel = 113;
			5127: Pixel = 110;
			5128: Pixel = 102;
			5129: Pixel = 92;
			5130: Pixel = 80;
			5131: Pixel = 75;
			5132: Pixel = 70;
			5133: Pixel = 61;
			5134: Pixel = 56;
			5135: Pixel = 51;
			5136: Pixel = 93;
			5137: Pixel = 139;
			5138: Pixel = 108;
			5139: Pixel = 126;
			5140: Pixel = 241;
			5141: Pixel = 248;
			5142: Pixel = 245;
			5143: Pixel = 248;
			5144: Pixel = 247;
			5145: Pixel = 208;
			5146: Pixel = 187;
			5147: Pixel = 187;
			5148: Pixel = 155;
			5149: Pixel = 182;
			5150: Pixel = 190;
			5151: Pixel = 160;
			5152: Pixel = 98;
			5153: Pixel = 66;
			5154: Pixel = 76;
			5155: Pixel = 77;
			5156: Pixel = 79;
			5157: Pixel = 84;
			5158: Pixel = 94;
			5159: Pixel = 115;
			5160: Pixel = 141;
			5161: Pixel = 159;
			5162: Pixel = 175;
			5163: Pixel = 189;
			5164: Pixel = 196;
			5165: Pixel = 200;
			5166: Pixel = 200;
			5167: Pixel = 156;
			5168: Pixel = 73;
			5169: Pixel = 70;
			5170: Pixel = 65;
			5171: Pixel = 49;
			5172: Pixel = 47;
			5173: Pixel = 53;
			5174: Pixel = 68;
			5175: Pixel = 55;
			5176: Pixel = 88;
			5177: Pixel = 70;
			5178: Pixel = 65;
			5179: Pixel = 63;
			5180: Pixel = 56;
			5181: Pixel = 56;
			5182: Pixel = 54;
			5183: Pixel = 57;
			5184: Pixel = 52;
			5185: Pixel = 65;
			5186: Pixel = 65;
			5187: Pixel = 68;
			5188: Pixel = 73;
			5189: Pixel = 56;
			5190: Pixel = 48;
			5191: Pixel = 93;
			5192: Pixel = 165;
			5193: Pixel = 231;
			5194: Pixel = 255;
			5195: Pixel = 229;
			5196: Pixel = 153;
			5197: Pixel = 87;
			5198: Pixel = 58;
			5199: Pixel = 65;
			5200: Pixel = 194;
			5201: Pixel = 184;
			5202: Pixel = 183;
			5203: Pixel = 185;
			5204: Pixel = 180;
			5205: Pixel = 167;
			5206: Pixel = 141;
			5207: Pixel = 157;
			5208: Pixel = 209;
			5209: Pixel = 218;
			5210: Pixel = 175;
			5211: Pixel = 142;
			5212: Pixel = 166;
			5213: Pixel = 189;
			5214: Pixel = 162;
			5215: Pixel = 166;
			5216: Pixel = 154;
			5217: Pixel = 137;
			5218: Pixel = 130;
			5219: Pixel = 113;
			5220: Pixel = 94;
			5221: Pixel = 100;
			5222: Pixel = 116;
			5223: Pixel = 106;
			5224: Pixel = 103;
			5225: Pixel = 110;
			5226: Pixel = 104;
			5227: Pixel = 96;
			5228: Pixel = 88;
			5229: Pixel = 74;
			5230: Pixel = 67;
			5231: Pixel = 65;
			5232: Pixel = 61;
			5233: Pixel = 61;
			5234: Pixel = 65;
			5235: Pixel = 59;
			5236: Pixel = 65;
			5237: Pixel = 115;
			5238: Pixel = 106;
			5239: Pixel = 101;
			5240: Pixel = 197;
			5241: Pixel = 254;
			5242: Pixel = 249;
			5243: Pixel = 241;
			5244: Pixel = 199;
			5245: Pixel = 184;
			5246: Pixel = 166;
			5247: Pixel = 126;
			5248: Pixel = 182;
			5249: Pixel = 175;
			5250: Pixel = 146;
			5251: Pixel = 156;
			5252: Pixel = 156;
			5253: Pixel = 84;
			5254: Pixel = 89;
			5255: Pixel = 107;
			5256: Pixel = 122;
			5257: Pixel = 133;
			5258: Pixel = 145;
			5259: Pixel = 159;
			5260: Pixel = 175;
			5261: Pixel = 186;
			5262: Pixel = 196;
			5263: Pixel = 203;
			5264: Pixel = 208;
			5265: Pixel = 202;
			5266: Pixel = 206;
			5267: Pixel = 201;
			5268: Pixel = 121;
			5269: Pixel = 66;
			5270: Pixel = 64;
			5271: Pixel = 48;
			5272: Pixel = 45;
			5273: Pixel = 53;
			5274: Pixel = 65;
			5275: Pixel = 54;
			5276: Pixel = 48;
			5277: Pixel = 53;
			5278: Pixel = 55;
			5279: Pixel = 56;
			5280: Pixel = 60;
			5281: Pixel = 65;
			5282: Pixel = 68;
			5283: Pixel = 67;
			5284: Pixel = 58;
			5285: Pixel = 66;
			5286: Pixel = 66;
			5287: Pixel = 64;
			5288: Pixel = 71;
			5289: Pixel = 115;
			5290: Pixel = 181;
			5291: Pixel = 245;
			5292: Pixel = 255;
			5293: Pixel = 228;
			5294: Pixel = 157;
			5295: Pixel = 82;
			5296: Pixel = 48;
			5297: Pixel = 54;
			5298: Pixel = 60;
			5299: Pixel = 56;
			5300: Pixel = 162;
			5301: Pixel = 155;
			5302: Pixel = 152;
			5303: Pixel = 153;
			5304: Pixel = 145;
			5305: Pixel = 140;
			5306: Pixel = 126;
			5307: Pixel = 179;
			5308: Pixel = 223;
			5309: Pixel = 179;
			5310: Pixel = 162;
			5311: Pixel = 160;
			5312: Pixel = 156;
			5313: Pixel = 151;
			5314: Pixel = 170;
			5315: Pixel = 174;
			5316: Pixel = 131;
			5317: Pixel = 122;
			5318: Pixel = 120;
			5319: Pixel = 115;
			5320: Pixel = 95;
			5321: Pixel = 111;
			5322: Pixel = 123;
			5323: Pixel = 108;
			5324: Pixel = 107;
			5325: Pixel = 101;
			5326: Pixel = 92;
			5327: Pixel = 82;
			5328: Pixel = 75;
			5329: Pixel = 76;
			5330: Pixel = 70;
			5331: Pixel = 68;
			5332: Pixel = 59;
			5333: Pixel = 56;
			5334: Pixel = 89;
			5335: Pixel = 62;
			5336: Pixel = 47;
			5337: Pixel = 100;
			5338: Pixel = 102;
			5339: Pixel = 98;
			5340: Pixel = 133;
			5341: Pixel = 255;
			5342: Pixel = 232;
			5343: Pixel = 188;
			5344: Pixel = 179;
			5345: Pixel = 154;
			5346: Pixel = 76;
			5347: Pixel = 158;
			5348: Pixel = 163;
			5349: Pixel = 143;
			5350: Pixel = 171;
			5351: Pixel = 192;
			5352: Pixel = 185;
			5353: Pixel = 130;
			5354: Pixel = 141;
			5355: Pixel = 160;
			5356: Pixel = 171;
			5357: Pixel = 182;
			5358: Pixel = 192;
			5359: Pixel = 196;
			5360: Pixel = 201;
			5361: Pixel = 202;
			5362: Pixel = 199;
			5363: Pixel = 202;
			5364: Pixel = 199;
			5365: Pixel = 207;
			5366: Pixel = 221;
			5367: Pixel = 218;
			5368: Pixel = 193;
			5369: Pixel = 107;
			5370: Pixel = 53;
			5371: Pixel = 47;
			5372: Pixel = 51;
			5373: Pixel = 53;
			5374: Pixel = 61;
			5375: Pixel = 53;
			5376: Pixel = 56;
			5377: Pixel = 60;
			5378: Pixel = 67;
			5379: Pixel = 70;
			5380: Pixel = 71;
			5381: Pixel = 72;
			5382: Pixel = 74;
			5383: Pixel = 72;
			5384: Pixel = 58;
			5385: Pixel = 62;
			5386: Pixel = 76;
			5387: Pixel = 125;
			5388: Pixel = 194;
			5389: Pixel = 250;
			5390: Pixel = 255;
			5391: Pixel = 221;
			5392: Pixel = 153;
			5393: Pixel = 84;
			5394: Pixel = 51;
			5395: Pixel = 47;
			5396: Pixel = 50;
			5397: Pixel = 50;
			5398: Pixel = 51;
			5399: Pixel = 47;
			5400: Pixel = 133;
			5401: Pixel = 134;
			5402: Pixel = 129;
			5403: Pixel = 127;
			5404: Pixel = 125;
			5405: Pixel = 127;
			5406: Pixel = 118;
			5407: Pixel = 141;
			5408: Pixel = 155;
			5409: Pixel = 169;
			5410: Pixel = 146;
			5411: Pixel = 144;
			5412: Pixel = 143;
			5413: Pixel = 134;
			5414: Pixel = 126;
			5415: Pixel = 163;
			5416: Pixel = 148;
			5417: Pixel = 119;
			5418: Pixel = 118;
			5419: Pixel = 118;
			5420: Pixel = 96;
			5421: Pixel = 113;
			5422: Pixel = 125;
			5423: Pixel = 122;
			5424: Pixel = 114;
			5425: Pixel = 106;
			5426: Pixel = 95;
			5427: Pixel = 84;
			5428: Pixel = 75;
			5429: Pixel = 70;
			5430: Pixel = 71;
			5431: Pixel = 69;
			5432: Pixel = 63;
			5433: Pixel = 71;
			5434: Pixel = 82;
			5435: Pixel = 57;
			5436: Pixel = 44;
			5437: Pixel = 72;
			5438: Pixel = 107;
			5439: Pixel = 104;
			5440: Pixel = 96;
			5441: Pixel = 191;
			5442: Pixel = 185;
			5443: Pixel = 182;
			5444: Pixel = 146;
			5445: Pixel = 108;
			5446: Pixel = 145;
			5447: Pixel = 119;
			5448: Pixel = 117;
			5449: Pixel = 159;
			5450: Pixel = 189;
			5451: Pixel = 194;
			5452: Pixel = 185;
			5453: Pixel = 163;
			5454: Pixel = 163;
			5455: Pixel = 188;
			5456: Pixel = 198;
			5457: Pixel = 190;
			5458: Pixel = 180;
			5459: Pixel = 176;
			5460: Pixel = 165;
			5461: Pixel = 150;
			5462: Pixel = 146;
			5463: Pixel = 146;
			5464: Pixel = 189;
			5465: Pixel = 224;
			5466: Pixel = 242;
			5467: Pixel = 217;
			5468: Pixel = 193;
			5469: Pixel = 166;
			5470: Pixel = 76;
			5471: Pixel = 44;
			5472: Pixel = 51;
			5473: Pixel = 56;
			5474: Pixel = 62;
			5475: Pixel = 56;
			5476: Pixel = 66;
			5477: Pixel = 67;
			5478: Pixel = 66;
			5479: Pixel = 70;
			5480: Pixel = 72;
			5481: Pixel = 75;
			5482: Pixel = 70;
			5483: Pixel = 61;
			5484: Pixel = 80;
			5485: Pixel = 144;
			5486: Pixel = 213;
			5487: Pixel = 255;
			5488: Pixel = 254;
			5489: Pixel = 208;
			5490: Pixel = 135;
			5491: Pixel = 89;
			5492: Pixel = 69;
			5493: Pixel = 48;
			5494: Pixel = 51;
			5495: Pixel = 54;
			5496: Pixel = 50;
			5497: Pixel = 47;
			5498: Pixel = 48;
			5499: Pixel = 45;
			5500: Pixel = 114;
			5501: Pixel = 114;
			5502: Pixel = 113;
			5503: Pixel = 114;
			5504: Pixel = 114;
			5505: Pixel = 110;
			5506: Pixel = 102;
			5507: Pixel = 100;
			5508: Pixel = 150;
			5509: Pixel = 171;
			5510: Pixel = 134;
			5511: Pixel = 136;
			5512: Pixel = 137;
			5513: Pixel = 128;
			5514: Pixel = 116;
			5515: Pixel = 155;
			5516: Pixel = 157;
			5517: Pixel = 137;
			5518: Pixel = 132;
			5519: Pixel = 116;
			5520: Pixel = 94;
			5521: Pixel = 114;
			5522: Pixel = 112;
			5523: Pixel = 117;
			5524: Pixel = 105;
			5525: Pixel = 104;
			5526: Pixel = 95;
			5527: Pixel = 81;
			5528: Pixel = 77;
			5529: Pixel = 77;
			5530: Pixel = 72;
			5531: Pixel = 65;
			5532: Pixel = 71;
			5533: Pixel = 82;
			5534: Pixel = 63;
			5535: Pixel = 49;
			5536: Pixel = 53;
			5537: Pixel = 56;
			5538: Pixel = 84;
			5539: Pixel = 95;
			5540: Pixel = 96;
			5541: Pixel = 122;
			5542: Pixel = 138;
			5543: Pixel = 157;
			5544: Pixel = 129;
			5545: Pixel = 117;
			5546: Pixel = 161;
			5547: Pixel = 151;
			5548: Pixel = 139;
			5549: Pixel = 164;
			5550: Pixel = 184;
			5551: Pixel = 187;
			5552: Pixel = 182;
			5553: Pixel = 177;
			5554: Pixel = 187;
			5555: Pixel = 202;
			5556: Pixel = 184;
			5557: Pixel = 153;
			5558: Pixel = 136;
			5559: Pixel = 128;
			5560: Pixel = 128;
			5561: Pixel = 126;
			5562: Pixel = 118;
			5563: Pixel = 136;
			5564: Pixel = 202;
			5565: Pixel = 224;
			5566: Pixel = 214;
			5567: Pixel = 202;
			5568: Pixel = 196;
			5569: Pixel = 165;
			5570: Pixel = 124;
			5571: Pixel = 53;
			5572: Pixel = 47;
			5573: Pixel = 57;
			5574: Pixel = 64;
			5575: Pixel = 59;
			5576: Pixel = 64;
			5577: Pixel = 62;
			5578: Pixel = 66;
			5579: Pixel = 69;
			5580: Pixel = 63;
			5581: Pixel = 64;
			5582: Pixel = 94;
			5583: Pixel = 155;
			5584: Pixel = 226;
			5585: Pixel = 255;
			5586: Pixel = 246;
			5587: Pixel = 192;
			5588: Pixel = 124;
			5589: Pixel = 76;
			5590: Pixel = 48;
			5591: Pixel = 65;
			5592: Pixel = 85;
			5593: Pixel = 67;
			5594: Pixel = 44;
			5595: Pixel = 42;
			5596: Pixel = 44;
			5597: Pixel = 45;
			5598: Pixel = 43;
			5599: Pixel = 38;
			5600: Pixel = 105;
			5601: Pixel = 103;
			5602: Pixel = 100;
			5603: Pixel = 96;
			5604: Pixel = 96;
			5605: Pixel = 107;
			5606: Pixel = 122;
			5607: Pixel = 150;
			5608: Pixel = 180;
			5609: Pixel = 165;
			5610: Pixel = 141;
			5611: Pixel = 134;
			5612: Pixel = 130;
			5613: Pixel = 124;
			5614: Pixel = 116;
			5615: Pixel = 155;
			5616: Pixel = 165;
			5617: Pixel = 153;
			5618: Pixel = 162;
			5619: Pixel = 127;
			5620: Pixel = 94;
			5621: Pixel = 137;
			5622: Pixel = 119;
			5623: Pixel = 110;
			5624: Pixel = 105;
			5625: Pixel = 98;
			5626: Pixel = 89;
			5627: Pixel = 83;
			5628: Pixel = 84;
			5629: Pixel = 100;
			5630: Pixel = 85;
			5631: Pixel = 63;
			5632: Pixel = 65;
			5633: Pixel = 70;
			5634: Pixel = 57;
			5635: Pixel = 52;
			5636: Pixel = 55;
			5637: Pixel = 57;
			5638: Pixel = 59;
			5639: Pixel = 69;
			5640: Pixel = 125;
			5641: Pixel = 147;
			5642: Pixel = 106;
			5643: Pixel = 137;
			5644: Pixel = 125;
			5645: Pixel = 125;
			5646: Pixel = 140;
			5647: Pixel = 163;
			5648: Pixel = 155;
			5649: Pixel = 153;
			5650: Pixel = 173;
			5651: Pixel = 183;
			5652: Pixel = 202;
			5653: Pixel = 223;
			5654: Pixel = 234;
			5655: Pixel = 231;
			5656: Pixel = 212;
			5657: Pixel = 157;
			5658: Pixel = 139;
			5659: Pixel = 132;
			5660: Pixel = 122;
			5661: Pixel = 121;
			5662: Pixel = 110;
			5663: Pixel = 130;
			5664: Pixel = 185;
			5665: Pixel = 191;
			5666: Pixel = 221;
			5667: Pixel = 200;
			5668: Pixel = 166;
			5669: Pixel = 167;
			5670: Pixel = 155;
			5671: Pixel = 71;
			5672: Pixel = 45;
			5673: Pixel = 63;
			5674: Pixel = 65;
			5675: Pixel = 60;
			5676: Pixel = 65;
			5677: Pixel = 64;
			5678: Pixel = 58;
			5679: Pixel = 64;
			5680: Pixel = 100;
			5681: Pixel = 171;
			5682: Pixel = 237;
			5683: Pixel = 255;
			5684: Pixel = 236;
			5685: Pixel = 175;
			5686: Pixel = 112;
			5687: Pixel = 70;
			5688: Pixel = 59;
			5689: Pixel = 62;
			5690: Pixel = 55;
			5691: Pixel = 72;
			5692: Pixel = 79;
			5693: Pixel = 67;
			5694: Pixel = 60;
			5695: Pixel = 43;
			5696: Pixel = 41;
			5697: Pixel = 44;
			5698: Pixel = 44;
			5699: Pixel = 42;
			5700: Pixel = 93;
			5701: Pixel = 93;
			5702: Pixel = 95;
			5703: Pixel = 110;
			5704: Pixel = 136;
			5705: Pixel = 161;
			5706: Pixel = 166;
			5707: Pixel = 181;
			5708: Pixel = 167;
			5709: Pixel = 163;
			5710: Pixel = 144;
			5711: Pixel = 135;
			5712: Pixel = 129;
			5713: Pixel = 126;
			5714: Pixel = 117;
			5715: Pixel = 152;
			5716: Pixel = 166;
			5717: Pixel = 158;
			5718: Pixel = 164;
			5719: Pixel = 133;
			5720: Pixel = 93;
			5721: Pixel = 129;
			5722: Pixel = 123;
			5723: Pixel = 116;
			5724: Pixel = 109;
			5725: Pixel = 105;
			5726: Pixel = 105;
			5727: Pixel = 88;
			5728: Pixel = 72;
			5729: Pixel = 69;
			5730: Pixel = 81;
			5731: Pixel = 70;
			5732: Pixel = 71;
			5733: Pixel = 67;
			5734: Pixel = 55;
			5735: Pixel = 52;
			5736: Pixel = 53;
			5737: Pixel = 54;
			5738: Pixel = 57;
			5739: Pixel = 68;
			5740: Pixel = 146;
			5741: Pixel = 166;
			5742: Pixel = 110;
			5743: Pixel = 119;
			5744: Pixel = 112;
			5745: Pixel = 118;
			5746: Pixel = 135;
			5747: Pixel = 155;
			5748: Pixel = 150;
			5749: Pixel = 143;
			5750: Pixel = 159;
			5751: Pixel = 202;
			5752: Pixel = 241;
			5753: Pixel = 249;
			5754: Pixel = 233;
			5755: Pixel = 221;
			5756: Pixel = 210;
			5757: Pixel = 151;
			5758: Pixel = 120;
			5759: Pixel = 129;
			5760: Pixel = 115;
			5761: Pixel = 114;
			5762: Pixel = 98;
			5763: Pixel = 120;
			5764: Pixel = 151;
			5765: Pixel = 186;
			5766: Pixel = 189;
			5767: Pixel = 156;
			5768: Pixel = 159;
			5769: Pixel = 152;
			5770: Pixel = 162;
			5771: Pixel = 84;
			5772: Pixel = 45;
			5773: Pixel = 68;
			5774: Pixel = 66;
			5775: Pixel = 62;
			5776: Pixel = 55;
			5777: Pixel = 61;
			5778: Pixel = 105;
			5779: Pixel = 182;
			5780: Pixel = 244;
			5781: Pixel = 255;
			5782: Pixel = 222;
			5783: Pixel = 158;
			5784: Pixel = 95;
			5785: Pixel = 62;
			5786: Pixel = 60;
			5787: Pixel = 64;
			5788: Pixel = 65;
			5789: Pixel = 59;
			5790: Pixel = 52;
			5791: Pixel = 73;
			5792: Pixel = 76;
			5793: Pixel = 61;
			5794: Pixel = 65;
			5795: Pixel = 62;
			5796: Pixel = 45;
			5797: Pixel = 39;
			5798: Pixel = 40;
			5799: Pixel = 43;
			5800: Pixel = 106;
			5801: Pixel = 127;
			5802: Pixel = 150;
			5803: Pixel = 155;
			5804: Pixel = 152;
			5805: Pixel = 149;
			5806: Pixel = 154;
			5807: Pixel = 160;
			5808: Pixel = 149;
			5809: Pixel = 164;
			5810: Pixel = 144;
			5811: Pixel = 139;
			5812: Pixel = 127;
			5813: Pixel = 138;
			5814: Pixel = 124;
			5815: Pixel = 147;
			5816: Pixel = 170;
			5817: Pixel = 176;
			5818: Pixel = 164;
			5819: Pixel = 139;
			5820: Pixel = 95;
			5821: Pixel = 130;
			5822: Pixel = 124;
			5823: Pixel = 118;
			5824: Pixel = 110;
			5825: Pixel = 110;
			5826: Pixel = 100;
			5827: Pixel = 85;
			5828: Pixel = 71;
			5829: Pixel = 69;
			5830: Pixel = 75;
			5831: Pixel = 80;
			5832: Pixel = 77;
			5833: Pixel = 63;
			5834: Pixel = 52;
			5835: Pixel = 49;
			5836: Pixel = 53;
			5837: Pixel = 55;
			5838: Pixel = 60;
			5839: Pixel = 89;
			5840: Pixel = 194;
			5841: Pixel = 183;
			5842: Pixel = 106;
			5843: Pixel = 93;
			5844: Pixel = 101;
			5845: Pixel = 110;
			5846: Pixel = 128;
			5847: Pixel = 148;
			5848: Pixel = 144;
			5849: Pixel = 142;
			5850: Pixel = 186;
			5851: Pixel = 243;
			5852: Pixel = 249;
			5853: Pixel = 247;
			5854: Pixel = 232;
			5855: Pixel = 217;
			5856: Pixel = 204;
			5857: Pixel = 176;
			5858: Pixel = 115;
			5859: Pixel = 118;
			5860: Pixel = 112;
			5861: Pixel = 111;
			5862: Pixel = 87;
			5863: Pixel = 104;
			5864: Pixel = 139;
			5865: Pixel = 176;
			5866: Pixel = 155;
			5867: Pixel = 161;
			5868: Pixel = 158;
			5869: Pixel = 153;
			5870: Pixel = 159;
			5871: Pixel = 84;
			5872: Pixel = 51;
			5873: Pixel = 68;
			5874: Pixel = 56;
			5875: Pixel = 63;
			5876: Pixel = 113;
			5877: Pixel = 191;
			5878: Pixel = 250;
			5879: Pixel = 255;
			5880: Pixel = 211;
			5881: Pixel = 144;
			5882: Pixel = 92;
			5883: Pixel = 65;
			5884: Pixel = 58;
			5885: Pixel = 62;
			5886: Pixel = 63;
			5887: Pixel = 60;
			5888: Pixel = 61;
			5889: Pixel = 54;
			5890: Pixel = 50;
			5891: Pixel = 75;
			5892: Pixel = 74;
			5893: Pixel = 58;
			5894: Pixel = 62;
			5895: Pixel = 64;
			5896: Pixel = 61;
			5897: Pixel = 44;
			5898: Pixel = 39;
			5899: Pixel = 41;
			5900: Pixel = 147;
			5901: Pixel = 150;
			5902: Pixel = 143;
			5903: Pixel = 133;
			5904: Pixel = 149;
			5905: Pixel = 144;
			5906: Pixel = 133;
			5907: Pixel = 154;
			5908: Pixel = 160;
			5909: Pixel = 159;
			5910: Pixel = 141;
			5911: Pixel = 141;
			5912: Pixel = 138;
			5913: Pixel = 135;
			5914: Pixel = 112;
			5915: Pixel = 165;
			5916: Pixel = 182;
			5917: Pixel = 186;
			5918: Pixel = 179;
			5919: Pixel = 163;
			5920: Pixel = 102;
			5921: Pixel = 154;
			5922: Pixel = 156;
			5923: Pixel = 130;
			5924: Pixel = 113;
			5925: Pixel = 109;
			5926: Pixel = 90;
			5927: Pixel = 78;
			5928: Pixel = 81;
			5929: Pixel = 71;
			5930: Pixel = 69;
			5931: Pixel = 73;
			5932: Pixel = 73;
			5933: Pixel = 54;
			5934: Pixel = 53;
			5935: Pixel = 47;
			5936: Pixel = 51;
			5937: Pixel = 54;
			5938: Pixel = 62;
			5939: Pixel = 121;
			5940: Pixel = 222;
			5941: Pixel = 187;
			5942: Pixel = 101;
			5943: Pixel = 91;
			5944: Pixel = 93;
			5945: Pixel = 99;
			5946: Pixel = 120;
			5947: Pixel = 141;
			5948: Pixel = 136;
			5949: Pixel = 154;
			5950: Pixel = 218;
			5951: Pixel = 250;
			5952: Pixel = 241;
			5953: Pixel = 220;
			5954: Pixel = 196;
			5955: Pixel = 168;
			5956: Pixel = 146;
			5957: Pixel = 149;
			5958: Pixel = 105;
			5959: Pixel = 102;
			5960: Pixel = 106;
			5961: Pixel = 106;
			5962: Pixel = 85;
			5963: Pixel = 87;
			5964: Pixel = 130;
			5965: Pixel = 157;
			5966: Pixel = 149;
			5967: Pixel = 150;
			5968: Pixel = 152;
			5969: Pixel = 160;
			5970: Pixel = 154;
			5971: Pixel = 60;
			5972: Pixel = 43;
			5973: Pixel = 73;
			5974: Pixel = 121;
			5975: Pixel = 201;
			5976: Pixel = 254;
			5977: Pixel = 248;
			5978: Pixel = 195;
			5979: Pixel = 129;
			5980: Pixel = 82;
			5981: Pixel = 67;
			5982: Pixel = 70;
			5983: Pixel = 68;
			5984: Pixel = 59;
			5985: Pixel = 59;
			5986: Pixel = 57;
			5987: Pixel = 55;
			5988: Pixel = 56;
			5989: Pixel = 49;
			5990: Pixel = 54;
			5991: Pixel = 77;
			5992: Pixel = 67;
			5993: Pixel = 50;
			5994: Pixel = 56;
			5995: Pixel = 60;
			5996: Pixel = 61;
			5997: Pixel = 63;
			5998: Pixel = 45;
			5999: Pixel = 37;
			6000: Pixel = 140;
			6001: Pixel = 132;
			6002: Pixel = 130;
			6003: Pixel = 135;
			6004: Pixel = 138;
			6005: Pixel = 144;
			6006: Pixel = 161;
			6007: Pixel = 138;
			6008: Pixel = 145;
			6009: Pixel = 165;
			6010: Pixel = 143;
			6011: Pixel = 141;
			6012: Pixel = 135;
			6013: Pixel = 132;
			6014: Pixel = 117;
			6015: Pixel = 146;
			6016: Pixel = 172;
			6017: Pixel = 155;
			6018: Pixel = 139;
			6019: Pixel = 154;
			6020: Pixel = 100;
			6021: Pixel = 143;
			6022: Pixel = 177;
			6023: Pixel = 162;
			6024: Pixel = 117;
			6025: Pixel = 105;
			6026: Pixel = 94;
			6027: Pixel = 107;
			6028: Pixel = 88;
			6029: Pixel = 71;
			6030: Pixel = 74;
			6031: Pixel = 88;
			6032: Pixel = 77;
			6033: Pixel = 49;
			6034: Pixel = 50;
			6035: Pixel = 46;
			6036: Pixel = 51;
			6037: Pixel = 56;
			6038: Pixel = 44;
			6039: Pixel = 145;
			6040: Pixel = 215;
			6041: Pixel = 171;
			6042: Pixel = 93;
			6043: Pixel = 97;
			6044: Pixel = 88;
			6045: Pixel = 90;
			6046: Pixel = 117;
			6047: Pixel = 135;
			6048: Pixel = 133;
			6049: Pixel = 173;
			6050: Pixel = 218;
			6051: Pixel = 229;
			6052: Pixel = 210;
			6053: Pixel = 179;
			6054: Pixel = 154;
			6055: Pixel = 133;
			6056: Pixel = 110;
			6057: Pixel = 124;
			6058: Pixel = 108;
			6059: Pixel = 95;
			6060: Pixel = 118;
			6061: Pixel = 103;
			6062: Pixel = 90;
			6063: Pixel = 78;
			6064: Pixel = 120;
			6065: Pixel = 157;
			6066: Pixel = 151;
			6067: Pixel = 150;
			6068: Pixel = 149;
			6069: Pixel = 158;
			6070: Pixel = 106;
			6071: Pixel = 61;
			6072: Pixel = 131;
			6073: Pixel = 213;
			6074: Pixel = 255;
			6075: Pixel = 240;
			6076: Pixel = 179;
			6077: Pixel = 114;
			6078: Pixel = 75;
			6079: Pixel = 65;
			6080: Pixel = 72;
			6081: Pixel = 74;
			6082: Pixel = 73;
			6083: Pixel = 64;
			6084: Pixel = 55;
			6085: Pixel = 57;
			6086: Pixel = 56;
			6087: Pixel = 53;
			6088: Pixel = 54;
			6089: Pixel = 47;
			6090: Pixel = 58;
			6091: Pixel = 81;
			6092: Pixel = 62;
			6093: Pixel = 49;
			6094: Pixel = 53;
			6095: Pixel = 59;
			6096: Pixel = 61;
			6097: Pixel = 66;
			6098: Pixel = 68;
			6099: Pixel = 48;
			6100: Pixel = 134;
			6101: Pixel = 126;
			6102: Pixel = 123;
			6103: Pixel = 119;
			6104: Pixel = 123;
			6105: Pixel = 141;
			6106: Pixel = 134;
			6107: Pixel = 138;
			6108: Pixel = 154;
			6109: Pixel = 171;
			6110: Pixel = 137;
			6111: Pixel = 134;
			6112: Pixel = 140;
			6113: Pixel = 130;
			6114: Pixel = 126;
			6115: Pixel = 133;
			6116: Pixel = 169;
			6117: Pixel = 155;
			6118: Pixel = 130;
			6119: Pixel = 142;
			6120: Pixel = 102;
			6121: Pixel = 121;
			6122: Pixel = 144;
			6123: Pixel = 120;
			6124: Pixel = 113;
			6125: Pixel = 107;
			6126: Pixel = 107;
			6127: Pixel = 107;
			6128: Pixel = 104;
			6129: Pixel = 100;
			6130: Pixel = 75;
			6131: Pixel = 83;
			6132: Pixel = 52;
			6133: Pixel = 49;
			6134: Pixel = 46;
			6135: Pixel = 46;
			6136: Pixel = 47;
			6137: Pixel = 51;
			6138: Pixel = 59;
			6139: Pixel = 155;
			6140: Pixel = 186;
			6141: Pixel = 142;
			6142: Pixel = 95;
			6143: Pixel = 100;
			6144: Pixel = 102;
			6145: Pixel = 87;
			6146: Pixel = 111;
			6147: Pixel = 128;
			6148: Pixel = 137;
			6149: Pixel = 170;
			6150: Pixel = 191;
			6151: Pixel = 205;
			6152: Pixel = 175;
			6153: Pixel = 159;
			6154: Pixel = 167;
			6155: Pixel = 172;
			6156: Pixel = 166;
			6157: Pixel = 119;
			6158: Pixel = 126;
			6159: Pixel = 184;
			6160: Pixel = 191;
			6161: Pixel = 100;
			6162: Pixel = 93;
			6163: Pixel = 71;
			6164: Pixel = 106;
			6165: Pixel = 157;
			6166: Pixel = 155;
			6167: Pixel = 151;
			6168: Pixel = 158;
			6169: Pixel = 150;
			6170: Pixel = 150;
			6171: Pixel = 217;
			6172: Pixel = 255;
			6173: Pixel = 229;
			6174: Pixel = 162;
			6175: Pixel = 100;
			6176: Pixel = 66;
			6177: Pixel = 62;
			6178: Pixel = 67;
			6179: Pixel = 68;
			6180: Pixel = 68;
			6181: Pixel = 69;
			6182: Pixel = 68;
			6183: Pixel = 61;
			6184: Pixel = 50;
			6185: Pixel = 54;
			6186: Pixel = 55;
			6187: Pixel = 51;
			6188: Pixel = 53;
			6189: Pixel = 46;
			6190: Pixel = 61;
			6191: Pixel = 79;
			6192: Pixel = 55;
			6193: Pixel = 47;
			6194: Pixel = 48;
			6195: Pixel = 49;
			6196: Pixel = 56;
			6197: Pixel = 62;
			6198: Pixel = 67;
			6199: Pixel = 65;
			6200: Pixel = 112;
			6201: Pixel = 134;
			6202: Pixel = 163;
			6203: Pixel = 129;
			6204: Pixel = 123;
			6205: Pixel = 130;
			6206: Pixel = 128;
			6207: Pixel = 157;
			6208: Pixel = 168;
			6209: Pixel = 169;
			6210: Pixel = 142;
			6211: Pixel = 137;
			6212: Pixel = 140;
			6213: Pixel = 136;
			6214: Pixel = 116;
			6215: Pixel = 111;
			6216: Pixel = 161;
			6217: Pixel = 151;
			6218: Pixel = 131;
			6219: Pixel = 139;
			6220: Pixel = 100;
			6221: Pixel = 96;
			6222: Pixel = 134;
			6223: Pixel = 119;
			6224: Pixel = 118;
			6225: Pixel = 125;
			6226: Pixel = 112;
			6227: Pixel = 85;
			6228: Pixel = 144;
			6229: Pixel = 145;
			6230: Pixel = 77;
			6231: Pixel = 67;
			6232: Pixel = 46;
			6233: Pixel = 48;
			6234: Pixel = 43;
			6235: Pixel = 48;
			6236: Pixel = 52;
			6237: Pixel = 50;
			6238: Pixel = 85;
			6239: Pixel = 160;
			6240: Pixel = 158;
			6241: Pixel = 124;
			6242: Pixel = 105;
			6243: Pixel = 104;
			6244: Pixel = 114;
			6245: Pixel = 108;
			6246: Pixel = 106;
			6247: Pixel = 123;
			6248: Pixel = 135;
			6249: Pixel = 149;
			6250: Pixel = 170;
			6251: Pixel = 174;
			6252: Pixel = 128;
			6253: Pixel = 165;
			6254: Pixel = 214;
			6255: Pixel = 223;
			6256: Pixel = 210;
			6257: Pixel = 179;
			6258: Pixel = 155;
			6259: Pixel = 214;
			6260: Pixel = 188;
			6261: Pixel = 103;
			6262: Pixel = 94;
			6263: Pixel = 74;
			6264: Pixel = 93;
			6265: Pixel = 134;
			6266: Pixel = 161;
			6267: Pixel = 152;
			6268: Pixel = 138;
			6269: Pixel = 169;
			6270: Pixel = 254;
			6271: Pixel = 214;
			6272: Pixel = 145;
			6273: Pixel = 92;
			6274: Pixel = 57;
			6275: Pixel = 60;
			6276: Pixel = 65;
			6277: Pixel = 65;
			6278: Pixel = 62;
			6279: Pixel = 63;
			6280: Pixel = 66;
			6281: Pixel = 66;
			6282: Pixel = 65;
			6283: Pixel = 58;
			6284: Pixel = 57;
			6285: Pixel = 58;
			6286: Pixel = 54;
			6287: Pixel = 51;
			6288: Pixel = 54;
			6289: Pixel = 46;
			6290: Pixel = 66;
			6291: Pixel = 79;
			6292: Pixel = 54;
			6293: Pixel = 46;
			6294: Pixel = 48;
			6295: Pixel = 47;
			6296: Pixel = 50;
			6297: Pixel = 57;
			6298: Pixel = 60;
			6299: Pixel = 62;
			6300: Pixel = 97;
			6301: Pixel = 108;
			6302: Pixel = 146;
			6303: Pixel = 156;
			6304: Pixel = 125;
			6305: Pixel = 122;
			6306: Pixel = 148;
			6307: Pixel = 171;
			6308: Pixel = 162;
			6309: Pixel = 171;
			6310: Pixel = 143;
			6311: Pixel = 135;
			6312: Pixel = 140;
			6313: Pixel = 139;
			6314: Pixel = 128;
			6315: Pixel = 118;
			6316: Pixel = 159;
			6317: Pixel = 157;
			6318: Pixel = 131;
			6319: Pixel = 135;
			6320: Pixel = 113;
			6321: Pixel = 88;
			6322: Pixel = 140;
			6323: Pixel = 140;
			6324: Pixel = 126;
			6325: Pixel = 120;
			6326: Pixel = 120;
			6327: Pixel = 101;
			6328: Pixel = 89;
			6329: Pixel = 93;
			6330: Pixel = 89;
			6331: Pixel = 53;
			6332: Pixel = 51;
			6333: Pixel = 46;
			6334: Pixel = 49;
			6335: Pixel = 47;
			6336: Pixel = 47;
			6337: Pixel = 48;
			6338: Pixel = 106;
			6339: Pixel = 161;
			6340: Pixel = 146;
			6341: Pixel = 116;
			6342: Pixel = 111;
			6343: Pixel = 110;
			6344: Pixel = 117;
			6345: Pixel = 124;
			6346: Pixel = 114;
			6347: Pixel = 116;
			6348: Pixel = 131;
			6349: Pixel = 134;
			6350: Pixel = 148;
			6351: Pixel = 127;
			6352: Pixel = 112;
			6353: Pixel = 185;
			6354: Pixel = 226;
			6355: Pixel = 214;
			6356: Pixel = 216;
			6357: Pixel = 222;
			6358: Pixel = 155;
			6359: Pixel = 160;
			6360: Pixel = 138;
			6361: Pixel = 98;
			6362: Pixel = 93;
			6363: Pixel = 85;
			6364: Pixel = 98;
			6365: Pixel = 94;
			6366: Pixel = 118;
			6367: Pixel = 125;
			6368: Pixel = 148;
			6369: Pixel = 163;
			6370: Pixel = 128;
			6371: Pixel = 65;
			6372: Pixel = 51;
			6373: Pixel = 67;
			6374: Pixel = 56;
			6375: Pixel = 57;
			6376: Pixel = 56;
			6377: Pixel = 58;
			6378: Pixel = 56;
			6379: Pixel = 57;
			6380: Pixel = 61;
			6381: Pixel = 60;
			6382: Pixel = 58;
			6383: Pixel = 52;
			6384: Pixel = 76;
			6385: Pixel = 64;
			6386: Pixel = 47;
			6387: Pixel = 49;
			6388: Pixel = 49;
			6389: Pixel = 39;
			6390: Pixel = 64;
			6391: Pixel = 79;
			6392: Pixel = 53;
			6393: Pixel = 49;
			6394: Pixel = 45;
			6395: Pixel = 44;
			6396: Pixel = 46;
			6397: Pixel = 46;
			6398: Pixel = 53;
			6399: Pixel = 56;
			6400: Pixel = 90;
			6401: Pixel = 91;
			6402: Pixel = 109;
			6403: Pixel = 133;
			6404: Pixel = 130;
			6405: Pixel = 134;
			6406: Pixel = 135;
			6407: Pixel = 145;
			6408: Pixel = 182;
			6409: Pixel = 162;
			6410: Pixel = 145;
			6411: Pixel = 138;
			6412: Pixel = 147;
			6413: Pixel = 146;
			6414: Pixel = 134;
			6415: Pixel = 109;
			6416: Pixel = 154;
			6417: Pixel = 148;
			6418: Pixel = 127;
			6419: Pixel = 142;
			6420: Pixel = 132;
			6421: Pixel = 81;
			6422: Pixel = 130;
			6423: Pixel = 129;
			6424: Pixel = 122;
			6425: Pixel = 132;
			6426: Pixel = 123;
			6427: Pixel = 127;
			6428: Pixel = 94;
			6429: Pixel = 92;
			6430: Pixel = 66;
			6431: Pixel = 49;
			6432: Pixel = 54;
			6433: Pixel = 50;
			6434: Pixel = 45;
			6435: Pixel = 87;
			6436: Pixel = 87;
			6437: Pixel = 49;
			6438: Pixel = 125;
			6439: Pixel = 157;
			6440: Pixel = 139;
			6441: Pixel = 115;
			6442: Pixel = 116;
			6443: Pixel = 115;
			6444: Pixel = 120;
			6445: Pixel = 127;
			6446: Pixel = 122;
			6447: Pixel = 117;
			6448: Pixel = 125;
			6449: Pixel = 123;
			6450: Pixel = 139;
			6451: Pixel = 116;
			6452: Pixel = 115;
			6453: Pixel = 202;
			6454: Pixel = 243;
			6455: Pixel = 220;
			6456: Pixel = 208;
			6457: Pixel = 199;
			6458: Pixel = 176;
			6459: Pixel = 129;
			6460: Pixel = 118;
			6461: Pixel = 95;
			6462: Pixel = 108;
			6463: Pixel = 108;
			6464: Pixel = 115;
			6465: Pixel = 114;
			6466: Pixel = 118;
			6467: Pixel = 149;
			6468: Pixel = 166;
			6469: Pixel = 138;
			6470: Pixel = 50;
			6471: Pixel = 44;
			6472: Pixel = 59;
			6473: Pixel = 67;
			6474: Pixel = 53;
			6475: Pixel = 53;
			6476: Pixel = 51;
			6477: Pixel = 55;
			6478: Pixel = 56;
			6479: Pixel = 53;
			6480: Pixel = 56;
			6481: Pixel = 57;
			6482: Pixel = 53;
			6483: Pixel = 51;
			6484: Pixel = 48;
			6485: Pixel = 51;
			6486: Pixel = 49;
			6487: Pixel = 49;
			6488: Pixel = 51;
			6489: Pixel = 40;
			6490: Pixel = 67;
			6491: Pixel = 76;
			6492: Pixel = 59;
			6493: Pixel = 60;
			6494: Pixel = 57;
			6495: Pixel = 48;
			6496: Pixel = 46;
			6497: Pixel = 48;
			6498: Pixel = 51;
			6499: Pixel = 53;
			6500: Pixel = 101;
			6501: Pixel = 111;
			6502: Pixel = 145;
			6503: Pixel = 138;
			6504: Pixel = 156;
			6505: Pixel = 171;
			6506: Pixel = 162;
			6507: Pixel = 165;
			6508: Pixel = 195;
			6509: Pixel = 152;
			6510: Pixel = 142;
			6511: Pixel = 149;
			6512: Pixel = 149;
			6513: Pixel = 138;
			6514: Pixel = 130;
			6515: Pixel = 99;
			6516: Pixel = 143;
			6517: Pixel = 137;
			6518: Pixel = 130;
			6519: Pixel = 152;
			6520: Pixel = 134;
			6521: Pixel = 76;
			6522: Pixel = 120;
			6523: Pixel = 127;
			6524: Pixel = 135;
			6525: Pixel = 161;
			6526: Pixel = 119;
			6527: Pixel = 121;
			6528: Pixel = 122;
			6529: Pixel = 77;
			6530: Pixel = 53;
			6531: Pixel = 65;
			6532: Pixel = 159;
			6533: Pixel = 142;
			6534: Pixel = 117;
			6535: Pixel = 173;
			6536: Pixel = 174;
			6537: Pixel = 80;
			6538: Pixel = 143;
			6539: Pixel = 154;
			6540: Pixel = 132;
			6541: Pixel = 118;
			6542: Pixel = 120;
			6543: Pixel = 118;
			6544: Pixel = 116;
			6545: Pixel = 124;
			6546: Pixel = 126;
			6547: Pixel = 121;
			6548: Pixel = 118;
			6549: Pixel = 111;
			6550: Pixel = 135;
			6551: Pixel = 108;
			6552: Pixel = 104;
			6553: Pixel = 163;
			6554: Pixel = 229;
			6555: Pixel = 202;
			6556: Pixel = 199;
			6557: Pixel = 193;
			6558: Pixel = 200;
			6559: Pixel = 131;
			6560: Pixel = 91;
			6561: Pixel = 91;
			6562: Pixel = 116;
			6563: Pixel = 115;
			6564: Pixel = 127;
			6565: Pixel = 133;
			6566: Pixel = 150;
			6567: Pixel = 166;
			6568: Pixel = 161;
			6569: Pixel = 129;
			6570: Pixel = 52;
			6571: Pixel = 44;
			6572: Pixel = 54;
			6573: Pixel = 59;
			6574: Pixel = 48;
			6575: Pixel = 50;
			6576: Pixel = 49;
			6577: Pixel = 52;
			6578: Pixel = 53;
			6579: Pixel = 50;
			6580: Pixel = 52;
			6581: Pixel = 52;
			6582: Pixel = 50;
			6583: Pixel = 46;
			6584: Pixel = 43;
			6585: Pixel = 47;
			6586: Pixel = 47;
			6587: Pixel = 49;
			6588: Pixel = 52;
			6589: Pixel = 41;
			6590: Pixel = 69;
			6591: Pixel = 76;
			6592: Pixel = 66;
			6593: Pixel = 68;
			6594: Pixel = 64;
			6595: Pixel = 54;
			6596: Pixel = 49;
			6597: Pixel = 48;
			6598: Pixel = 50;
			6599: Pixel = 49;
			6600: Pixel = 124;
			6601: Pixel = 124;
			6602: Pixel = 159;
			6603: Pixel = 150;
			6604: Pixel = 153;
			6605: Pixel = 193;
			6606: Pixel = 166;
			6607: Pixel = 186;
			6608: Pixel = 196;
			6609: Pixel = 179;
			6610: Pixel = 157;
			6611: Pixel = 149;
			6612: Pixel = 140;
			6613: Pixel = 141;
			6614: Pixel = 143;
			6615: Pixel = 99;
			6616: Pixel = 147;
			6617: Pixel = 140;
			6618: Pixel = 134;
			6619: Pixel = 153;
			6620: Pixel = 145;
			6621: Pixel = 82;
			6622: Pixel = 121;
			6623: Pixel = 137;
			6624: Pixel = 161;
			6625: Pixel = 139;
			6626: Pixel = 143;
			6627: Pixel = 144;
			6628: Pixel = 77;
			6629: Pixel = 56;
			6630: Pixel = 119;
			6631: Pixel = 219;
			6632: Pixel = 219;
			6633: Pixel = 181;
			6634: Pixel = 200;
			6635: Pixel = 200;
			6636: Pixel = 195;
			6637: Pixel = 133;
			6638: Pixel = 178;
			6639: Pixel = 157;
			6640: Pixel = 126;
			6641: Pixel = 119;
			6642: Pixel = 123;
			6643: Pixel = 122;
			6644: Pixel = 119;
			6645: Pixel = 125;
			6646: Pixel = 124;
			6647: Pixel = 127;
			6648: Pixel = 113;
			6649: Pixel = 100;
			6650: Pixel = 128;
			6651: Pixel = 109;
			6652: Pixel = 99;
			6653: Pixel = 94;
			6654: Pixel = 188;
			6655: Pixel = 209;
			6656: Pixel = 194;
			6657: Pixel = 196;
			6658: Pixel = 194;
			6659: Pixel = 177;
			6660: Pixel = 197;
			6661: Pixel = 86;
			6662: Pixel = 88;
			6663: Pixel = 106;
			6664: Pixel = 135;
			6665: Pixel = 137;
			6666: Pixel = 157;
			6667: Pixel = 161;
			6668: Pixel = 155;
			6669: Pixel = 103;
			6670: Pixel = 44;
			6671: Pixel = 41;
			6672: Pixel = 54;
			6673: Pixel = 52;
			6674: Pixel = 44;
			6675: Pixel = 47;
			6676: Pixel = 47;
			6677: Pixel = 49;
			6678: Pixel = 49;
			6679: Pixel = 48;
			6680: Pixel = 50;
			6681: Pixel = 49;
			6682: Pixel = 48;
			6683: Pixel = 47;
			6684: Pixel = 43;
			6685: Pixel = 45;
			6686: Pixel = 44;
			6687: Pixel = 46;
			6688: Pixel = 51;
			6689: Pixel = 43;
			6690: Pixel = 71;
			6691: Pixel = 79;
			6692: Pixel = 70;
			6693: Pixel = 76;
			6694: Pixel = 72;
			6695: Pixel = 63;
			6696: Pixel = 54;
			6697: Pixel = 51;
			6698: Pixel = 49;
			6699: Pixel = 48;
			6700: Pixel = 143;
			6701: Pixel = 146;
			6702: Pixel = 143;
			6703: Pixel = 163;
			6704: Pixel = 160;
			6705: Pixel = 154;
			6706: Pixel = 175;
			6707: Pixel = 217;
			6708: Pixel = 210;
			6709: Pixel = 190;
			6710: Pixel = 162;
			6711: Pixel = 144;
			6712: Pixel = 149;
			6713: Pixel = 153;
			6714: Pixel = 151;
			6715: Pixel = 107;
			6716: Pixel = 144;
			6717: Pixel = 141;
			6718: Pixel = 133;
			6719: Pixel = 146;
			6720: Pixel = 157;
			6721: Pixel = 82;
			6722: Pixel = 128;
			6723: Pixel = 159;
			6724: Pixel = 164;
			6725: Pixel = 144;
			6726: Pixel = 125;
			6727: Pixel = 85;
			6728: Pixel = 70;
			6729: Pixel = 56;
			6730: Pixel = 130;
			6731: Pixel = 185;
			6732: Pixel = 164;
			6733: Pixel = 179;
			6734: Pixel = 212;
			6735: Pixel = 210;
			6736: Pixel = 213;
			6737: Pixel = 175;
			6738: Pixel = 201;
			6739: Pixel = 155;
			6740: Pixel = 118;
			6741: Pixel = 122;
			6742: Pixel = 122;
			6743: Pixel = 124;
			6744: Pixel = 121;
			6745: Pixel = 123;
			6746: Pixel = 127;
			6747: Pixel = 113;
			6748: Pixel = 105;
			6749: Pixel = 99;
			6750: Pixel = 119;
			6751: Pixel = 112;
			6752: Pixel = 93;
			6753: Pixel = 84;
			6754: Pixel = 130;
			6755: Pixel = 213;
			6756: Pixel = 193;
			6757: Pixel = 198;
			6758: Pixel = 201;
			6759: Pixel = 227;
			6760: Pixel = 212;
			6761: Pixel = 92;
			6762: Pixel = 65;
			6763: Pixel = 98;
			6764: Pixel = 139;
			6765: Pixel = 144;
			6766: Pixel = 153;
			6767: Pixel = 144;
			6768: Pixel = 128;
			6769: Pixel = 65;
			6770: Pixel = 45;
			6771: Pixel = 38;
			6772: Pixel = 50;
			6773: Pixel = 48;
			6774: Pixel = 43;
			6775: Pixel = 44;
			6776: Pixel = 44;
			6777: Pixel = 46;
			6778: Pixel = 46;
			6779: Pixel = 45;
			6780: Pixel = 48;
			6781: Pixel = 48;
			6782: Pixel = 45;
			6783: Pixel = 44;
			6784: Pixel = 39;
			6785: Pixel = 42;
			6786: Pixel = 40;
			6787: Pixel = 41;
			6788: Pixel = 43;
			6789: Pixel = 41;
			6790: Pixel = 74;
			6791: Pixel = 74;
			6792: Pixel = 74;
			6793: Pixel = 80;
			6794: Pixel = 76;
			6795: Pixel = 68;
			6796: Pixel = 61;
			6797: Pixel = 54;
			6798: Pixel = 54;
			6799: Pixel = 48;
			6800: Pixel = 169;
			6801: Pixel = 163;
			6802: Pixel = 183;
			6803: Pixel = 201;
			6804: Pixel = 191;
			6805: Pixel = 187;
			6806: Pixel = 173;
			6807: Pixel = 213;
			6808: Pixel = 243;
			6809: Pixel = 197;
			6810: Pixel = 152;
			6811: Pixel = 163;
			6812: Pixel = 164;
			6813: Pixel = 164;
			6814: Pixel = 177;
			6815: Pixel = 153;
			6816: Pixel = 125;
			6817: Pixel = 159;
			6818: Pixel = 145;
			6819: Pixel = 161;
			6820: Pixel = 185;
			6821: Pixel = 114;
			6822: Pixel = 133;
			6823: Pixel = 160;
			6824: Pixel = 120;
			6825: Pixel = 99;
			6826: Pixel = 66;
			6827: Pixel = 68;
			6828: Pixel = 73;
			6829: Pixel = 65;
			6830: Pixel = 76;
			6831: Pixel = 88;
			6832: Pixel = 129;
			6833: Pixel = 152;
			6834: Pixel = 183;
			6835: Pixel = 195;
			6836: Pixel = 157;
			6837: Pixel = 164;
			6838: Pixel = 176;
			6839: Pixel = 138;
			6840: Pixel = 120;
			6841: Pixel = 124;
			6842: Pixel = 124;
			6843: Pixel = 127;
			6844: Pixel = 125;
			6845: Pixel = 126;
			6846: Pixel = 131;
			6847: Pixel = 89;
			6848: Pixel = 76;
			6849: Pixel = 103;
			6850: Pixel = 112;
			6851: Pixel = 116;
			6852: Pixel = 97;
			6853: Pixel = 87;
			6854: Pixel = 87;
			6855: Pixel = 204;
			6856: Pixel = 218;
			6857: Pixel = 219;
			6858: Pixel = 208;
			6859: Pixel = 199;
			6860: Pixel = 106;
			6861: Pixel = 74;
			6862: Pixel = 88;
			6863: Pixel = 95;
			6864: Pixel = 129;
			6865: Pixel = 131;
			6866: Pixel = 130;
			6867: Pixel = 126;
			6868: Pixel = 79;
			6869: Pixel = 51;
			6870: Pixel = 49;
			6871: Pixel = 38;
			6872: Pixel = 46;
			6873: Pixel = 46;
			6874: Pixel = 45;
			6875: Pixel = 43;
			6876: Pixel = 44;
			6877: Pixel = 46;
			6878: Pixel = 48;
			6879: Pixel = 48;
			6880: Pixel = 47;
			6881: Pixel = 47;
			6882: Pixel = 47;
			6883: Pixel = 43;
			6884: Pixel = 40;
			6885: Pixel = 41;
			6886: Pixel = 41;
			6887: Pixel = 43;
			6888: Pixel = 36;
			6889: Pixel = 42;
			6890: Pixel = 78;
			6891: Pixel = 99;
			6892: Pixel = 78;
			6893: Pixel = 81;
			6894: Pixel = 79;
			6895: Pixel = 74;
			6896: Pixel = 68;
			6897: Pixel = 60;
			6898: Pixel = 56;
			6899: Pixel = 51;
			6900: Pixel = 189;
			6901: Pixel = 196;
			6902: Pixel = 197;
			6903: Pixel = 194;
			6904: Pixel = 211;
			6905: Pixel = 233;
			6906: Pixel = 223;
			6907: Pixel = 199;
			6908: Pixel = 237;
			6909: Pixel = 197;
			6910: Pixel = 164;
			6911: Pixel = 176;
			6912: Pixel = 174;
			6913: Pixel = 188;
			6914: Pixel = 184;
			6915: Pixel = 116;
			6916: Pixel = 132;
			6917: Pixel = 179;
			6918: Pixel = 172;
			6919: Pixel = 149;
			6920: Pixel = 119;
			6921: Pixel = 81;
			6922: Pixel = 88;
			6923: Pixel = 78;
			6924: Pixel = 66;
			6925: Pixel = 65;
			6926: Pixel = 70;
			6927: Pixel = 69;
			6928: Pixel = 68;
			6929: Pixel = 66;
			6930: Pixel = 67;
			6931: Pixel = 83;
			6932: Pixel = 106;
			6933: Pixel = 105;
			6934: Pixel = 96;
			6935: Pixel = 117;
			6936: Pixel = 127;
			6937: Pixel = 135;
			6938: Pixel = 140;
			6939: Pixel = 130;
			6940: Pixel = 124;
			6941: Pixel = 125;
			6942: Pixel = 124;
			6943: Pixel = 125;
			6944: Pixel = 125;
			6945: Pixel = 127;
			6946: Pixel = 121;
			6947: Pixel = 100;
			6948: Pixel = 84;
			6949: Pixel = 87;
			6950: Pixel = 94;
			6951: Pixel = 99;
			6952: Pixel = 99;
			6953: Pixel = 98;
			6954: Pixel = 82;
			6955: Pixel = 170;
			6956: Pixel = 228;
			6957: Pixel = 175;
			6958: Pixel = 144;
			6959: Pixel = 144;
			6960: Pixel = 107;
			6961: Pixel = 72;
			6962: Pixel = 85;
			6963: Pixel = 96;
			6964: Pixel = 116;
			6965: Pixel = 118;
			6966: Pixel = 124;
			6967: Pixel = 110;
			6968: Pixel = 50;
			6969: Pixel = 51;
			6970: Pixel = 46;
			6971: Pixel = 37;
			6972: Pixel = 43;
			6973: Pixel = 47;
			6974: Pixel = 45;
			6975: Pixel = 45;
			6976: Pixel = 44;
			6977: Pixel = 45;
			6978: Pixel = 45;
			6979: Pixel = 45;
			6980: Pixel = 44;
			6981: Pixel = 44;
			6982: Pixel = 43;
			6983: Pixel = 39;
			6984: Pixel = 41;
			6985: Pixel = 40;
			6986: Pixel = 39;
			6987: Pixel = 38;
			6988: Pixel = 59;
			6989: Pixel = 59;
			6990: Pixel = 93;
			6991: Pixel = 86;
			6992: Pixel = 74;
			6993: Pixel = 81;
			6994: Pixel = 79;
			6995: Pixel = 75;
			6996: Pixel = 70;
			6997: Pixel = 65;
			6998: Pixel = 60;
			6999: Pixel = 52;
			7000: Pixel = 225;
			7001: Pixel = 225;
			7002: Pixel = 206;
			7003: Pixel = 203;
			7004: Pixel = 216;
			7005: Pixel = 231;
			7006: Pixel = 220;
			7007: Pixel = 205;
			7008: Pixel = 195;
			7009: Pixel = 199;
			7010: Pixel = 194;
			7011: Pixel = 163;
			7012: Pixel = 143;
			7013: Pixel = 111;
			7014: Pixel = 77;
			7015: Pixel = 63;
			7016: Pixel = 130;
			7017: Pixel = 119;
			7018: Pixel = 90;
			7019: Pixel = 72;
			7020: Pixel = 66;
			7021: Pixel = 66;
			7022: Pixel = 64;
			7023: Pixel = 72;
			7024: Pixel = 71;
			7025: Pixel = 66;
			7026: Pixel = 67;
			7027: Pixel = 68;
			7028: Pixel = 66;
			7029: Pixel = 70;
			7030: Pixel = 69;
			7031: Pixel = 70;
			7032: Pixel = 55;
			7033: Pixel = 73;
			7034: Pixel = 164;
			7035: Pixel = 130;
			7036: Pixel = 130;
			7037: Pixel = 145;
			7038: Pixel = 148;
			7039: Pixel = 130;
			7040: Pixel = 124;
			7041: Pixel = 126;
			7042: Pixel = 125;
			7043: Pixel = 124;
			7044: Pixel = 125;
			7045: Pixel = 124;
			7046: Pixel = 128;
			7047: Pixel = 122;
			7048: Pixel = 102;
			7049: Pixel = 104;
			7050: Pixel = 144;
			7051: Pixel = 183;
			7052: Pixel = 151;
			7053: Pixel = 115;
			7054: Pixel = 97;
			7055: Pixel = 114;
			7056: Pixel = 146;
			7057: Pixel = 127;
			7058: Pixel = 97;
			7059: Pixel = 148;
			7060: Pixel = 117;
			7061: Pixel = 77;
			7062: Pixel = 80;
			7063: Pixel = 96;
			7064: Pixel = 118;
			7065: Pixel = 120;
			7066: Pixel = 140;
			7067: Pixel = 119;
			7068: Pixel = 47;
			7069: Pixel = 51;
			7070: Pixel = 48;
			7071: Pixel = 39;
			7072: Pixel = 45;
			7073: Pixel = 45;
			7074: Pixel = 44;
			7075: Pixel = 45;
			7076: Pixel = 44;
			7077: Pixel = 45;
			7078: Pixel = 45;
			7079: Pixel = 44;
			7080: Pixel = 46;
			7081: Pixel = 43;
			7082: Pixel = 43;
			7083: Pixel = 40;
			7084: Pixel = 39;
			7085: Pixel = 41;
			7086: Pixel = 39;
			7087: Pixel = 37;
			7088: Pixel = 72;
			7089: Pixel = 81;
			7090: Pixel = 96;
			7091: Pixel = 57;
			7092: Pixel = 72;
			7093: Pixel = 82;
			7094: Pixel = 78;
			7095: Pixel = 76;
			7096: Pixel = 71;
			7097: Pixel = 72;
			7098: Pixel = 68;
			7099: Pixel = 62;
			7100: Pixel = 188;
			7101: Pixel = 248;
			7102: Pixel = 219;
			7103: Pixel = 228;
			7104: Pixel = 204;
			7105: Pixel = 204;
			7106: Pixel = 174;
			7107: Pixel = 149;
			7108: Pixel = 103;
			7109: Pixel = 126;
			7110: Pixel = 118;
			7111: Pixel = 85;
			7112: Pixel = 73;
			7113: Pixel = 67;
			7114: Pixel = 70;
			7115: Pixel = 71;
			7116: Pixel = 67;
			7117: Pixel = 59;
			7118: Pixel = 61;
			7119: Pixel = 65;
			7120: Pixel = 64;
			7121: Pixel = 63;
			7122: Pixel = 65;
			7123: Pixel = 68;
			7124: Pixel = 62;
			7125: Pixel = 58;
			7126: Pixel = 57;
			7127: Pixel = 66;
			7128: Pixel = 73;
			7129: Pixel = 77;
			7130: Pixel = 76;
			7131: Pixel = 75;
			7132: Pixel = 56;
			7133: Pixel = 98;
			7134: Pixel = 205;
			7135: Pixel = 143;
			7136: Pixel = 135;
			7137: Pixel = 163;
			7138: Pixel = 156;
			7139: Pixel = 127;
			7140: Pixel = 127;
			7141: Pixel = 126;
			7142: Pixel = 127;
			7143: Pixel = 124;
			7144: Pixel = 124;
			7145: Pixel = 131;
			7146: Pixel = 172;
			7147: Pixel = 175;
			7148: Pixel = 154;
			7149: Pixel = 168;
			7150: Pixel = 195;
			7151: Pixel = 169;
			7152: Pixel = 122;
			7153: Pixel = 81;
			7154: Pixel = 64;
			7155: Pixel = 97;
			7156: Pixel = 145;
			7157: Pixel = 142;
			7158: Pixel = 164;
			7159: Pixel = 154;
			7160: Pixel = 123;
			7161: Pixel = 80;
			7162: Pixel = 88;
			7163: Pixel = 108;
			7164: Pixel = 145;
			7165: Pixel = 149;
			7166: Pixel = 156;
			7167: Pixel = 113;
			7168: Pixel = 45;
			7169: Pixel = 48;
			7170: Pixel = 48;
			7171: Pixel = 39;
			7172: Pixel = 46;
			7173: Pixel = 42;
			7174: Pixel = 42;
			7175: Pixel = 42;
			7176: Pixel = 41;
			7177: Pixel = 41;
			7178: Pixel = 42;
			7179: Pixel = 42;
			7180: Pixel = 43;
			7181: Pixel = 44;
			7182: Pixel = 38;
			7183: Pixel = 70;
			7184: Pixel = 52;
			7185: Pixel = 33;
			7186: Pixel = 37;
			7187: Pixel = 37;
			7188: Pixel = 29;
			7189: Pixel = 54;
			7190: Pixel = 74;
			7191: Pixel = 44;
			7192: Pixel = 56;
			7193: Pixel = 75;
			7194: Pixel = 77;
			7195: Pixel = 75;
			7196: Pixel = 72;
			7197: Pixel = 72;
			7198: Pixel = 71;
			7199: Pixel = 69;
			7200: Pixel = 103;
			7201: Pixel = 211;
			7202: Pixel = 201;
			7203: Pixel = 199;
			7204: Pixel = 172;
			7205: Pixel = 123;
			7206: Pixel = 89;
			7207: Pixel = 77;
			7208: Pixel = 78;
			7209: Pixel = 64;
			7210: Pixel = 66;
			7211: Pixel = 70;
			7212: Pixel = 81;
			7213: Pixel = 77;
			7214: Pixel = 72;
			7215: Pixel = 67;
			7216: Pixel = 62;
			7217: Pixel = 65;
			7218: Pixel = 65;
			7219: Pixel = 62;
			7220: Pixel = 60;
			7221: Pixel = 63;
			7222: Pixel = 63;
			7223: Pixel = 59;
			7224: Pixel = 55;
			7225: Pixel = 49;
			7226: Pixel = 54;
			7227: Pixel = 67;
			7228: Pixel = 78;
			7229: Pixel = 80;
			7230: Pixel = 73;
			7231: Pixel = 76;
			7232: Pixel = 56;
			7233: Pixel = 126;
			7234: Pixel = 183;
			7235: Pixel = 145;
			7236: Pixel = 160;
			7237: Pixel = 158;
			7238: Pixel = 134;
			7239: Pixel = 129;
			7240: Pixel = 126;
			7241: Pixel = 128;
			7242: Pixel = 128;
			7243: Pixel = 129;
			7244: Pixel = 118;
			7245: Pixel = 169;
			7246: Pixel = 227;
			7247: Pixel = 224;
			7248: Pixel = 219;
			7249: Pixel = 199;
			7250: Pixel = 158;
			7251: Pixel = 177;
			7252: Pixel = 137;
			7253: Pixel = 130;
			7254: Pixel = 122;
			7255: Pixel = 107;
			7256: Pixel = 134;
			7257: Pixel = 152;
			7258: Pixel = 153;
			7259: Pixel = 144;
			7260: Pixel = 91;
			7261: Pixel = 77;
			7262: Pixel = 89;
			7263: Pixel = 119;
			7264: Pixel = 155;
			7265: Pixel = 155;
			7266: Pixel = 157;
			7267: Pixel = 115;
			7268: Pixel = 46;
			7269: Pixel = 49;
			7270: Pixel = 47;
			7271: Pixel = 41;
			7272: Pixel = 49;
			7273: Pixel = 46;
			7274: Pixel = 44;
			7275: Pixel = 43;
			7276: Pixel = 43;
			7277: Pixel = 43;
			7278: Pixel = 41;
			7279: Pixel = 41;
			7280: Pixel = 43;
			7281: Pixel = 45;
			7282: Pixel = 44;
			7283: Pixel = 53;
			7284: Pixel = 44;
			7285: Pixel = 37;
			7286: Pixel = 38;
			7287: Pixel = 37;
			7288: Pixel = 33;
			7289: Pixel = 65;
			7290: Pixel = 79;
			7291: Pixel = 44;
			7292: Pixel = 48;
			7293: Pixel = 62;
			7294: Pixel = 80;
			7295: Pixel = 79;
			7296: Pixel = 76;
			7297: Pixel = 75;
			7298: Pixel = 72;
			7299: Pixel = 73;
			7300: Pixel = 74;
			7301: Pixel = 115;
			7302: Pixel = 115;
			7303: Pixel = 89;
			7304: Pixel = 74;
			7305: Pixel = 71;
			7306: Pixel = 73;
			7307: Pixel = 79;
			7308: Pixel = 71;
			7309: Pixel = 65;
			7310: Pixel = 70;
			7311: Pixel = 65;
			7312: Pixel = 76;
			7313: Pixel = 71;
			7314: Pixel = 66;
			7315: Pixel = 62;
			7316: Pixel = 60;
			7317: Pixel = 60;
			7318: Pixel = 62;
			7319: Pixel = 61;
			7320: Pixel = 61;
			7321: Pixel = 65;
			7322: Pixel = 60;
			7323: Pixel = 52;
			7324: Pixel = 55;
			7325: Pixel = 51;
			7326: Pixel = 57;
			7327: Pixel = 70;
			7328: Pixel = 72;
			7329: Pixel = 92;
			7330: Pixel = 132;
			7331: Pixel = 108;
			7332: Pixel = 85;
			7333: Pixel = 166;
			7334: Pixel = 183;
			7335: Pixel = 169;
			7336: Pixel = 197;
			7337: Pixel = 163;
			7338: Pixel = 128;
			7339: Pixel = 130;
			7340: Pixel = 129;
			7341: Pixel = 131;
			7342: Pixel = 130;
			7343: Pixel = 125;
			7344: Pixel = 124;
			7345: Pixel = 141;
			7346: Pixel = 159;
			7347: Pixel = 176;
			7348: Pixel = 185;
			7349: Pixel = 190;
			7350: Pixel = 126;
			7351: Pixel = 204;
			7352: Pixel = 238;
			7353: Pixel = 227;
			7354: Pixel = 228;
			7355: Pixel = 202;
			7356: Pixel = 139;
			7357: Pixel = 157;
			7358: Pixel = 172;
			7359: Pixel = 165;
			7360: Pixel = 133;
			7361: Pixel = 115;
			7362: Pixel = 80;
			7363: Pixel = 121;
			7364: Pixel = 155;
			7365: Pixel = 155;
			7366: Pixel = 158;
			7367: Pixel = 116;
			7368: Pixel = 41;
			7369: Pixel = 45;
			7370: Pixel = 41;
			7371: Pixel = 37;
			7372: Pixel = 41;
			7373: Pixel = 41;
			7374: Pixel = 43;
			7375: Pixel = 44;
			7376: Pixel = 45;
			7377: Pixel = 46;
			7378: Pixel = 42;
			7379: Pixel = 41;
			7380: Pixel = 45;
			7381: Pixel = 43;
			7382: Pixel = 45;
			7383: Pixel = 39;
			7384: Pixel = 38;
			7385: Pixel = 40;
			7386: Pixel = 36;
			7387: Pixel = 37;
			7388: Pixel = 34;
			7389: Pixel = 71;
			7390: Pixel = 76;
			7391: Pixel = 41;
			7392: Pixel = 45;
			7393: Pixel = 51;
			7394: Pixel = 71;
			7395: Pixel = 85;
			7396: Pixel = 79;
			7397: Pixel = 74;
			7398: Pixel = 72;
			7399: Pixel = 68;
			7400: Pixel = 69;
			7401: Pixel = 63;
			7402: Pixel = 60;
			7403: Pixel = 66;
			7404: Pixel = 71;
			7405: Pixel = 72;
			7406: Pixel = 73;
			7407: Pixel = 73;
			7408: Pixel = 71;
			7409: Pixel = 69;
			7410: Pixel = 67;
			7411: Pixel = 66;
			7412: Pixel = 63;
			7413: Pixel = 65;
			7414: Pixel = 63;
			7415: Pixel = 62;
			7416: Pixel = 58;
			7417: Pixel = 58;
			7418: Pixel = 62;
			7419: Pixel = 61;
			7420: Pixel = 61;
			7421: Pixel = 64;
			7422: Pixel = 62;
			7423: Pixel = 53;
			7424: Pixel = 56;
			7425: Pixel = 54;
			7426: Pixel = 66;
			7427: Pixel = 62;
			7428: Pixel = 99;
			7429: Pixel = 181;
			7430: Pixel = 231;
			7431: Pixel = 230;
			7432: Pixel = 217;
			7433: Pixel = 213;
			7434: Pixel = 208;
			7435: Pixel = 183;
			7436: Pixel = 219;
			7437: Pixel = 178;
			7438: Pixel = 132;
			7439: Pixel = 132;
			7440: Pixel = 132;
			7441: Pixel = 133;
			7442: Pixel = 127;
			7443: Pixel = 123;
			7444: Pixel = 121;
			7445: Pixel = 123;
			7446: Pixel = 128;
			7447: Pixel = 130;
			7448: Pixel = 164;
			7449: Pixel = 174;
			7450: Pixel = 79;
			7451: Pixel = 139;
			7452: Pixel = 171;
			7453: Pixel = 179;
			7454: Pixel = 197;
			7455: Pixel = 214;
			7456: Pixel = 195;
			7457: Pixel = 211;
			7458: Pixel = 230;
			7459: Pixel = 224;
			7460: Pixel = 233;
			7461: Pixel = 184;
			7462: Pixel = 73;
			7463: Pixel = 124;
			7464: Pixel = 155;
			7465: Pixel = 157;
			7466: Pixel = 153;
			7467: Pixel = 131;
			7468: Pixel = 104;
			7469: Pixel = 89;
			7470: Pixel = 73;
			7471: Pixel = 92;
			7472: Pixel = 98;
			7473: Pixel = 76;
			7474: Pixel = 56;
			7475: Pixel = 44;
			7476: Pixel = 41;
			7477: Pixel = 41;
			7478: Pixel = 40;
			7479: Pixel = 41;
			7480: Pixel = 43;
			7481: Pixel = 45;
			7482: Pixel = 45;
			7483: Pixel = 41;
			7484: Pixel = 42;
			7485: Pixel = 42;
			7486: Pixel = 41;
			7487: Pixel = 40;
			7488: Pixel = 38;
			7489: Pixel = 75;
			7490: Pixel = 73;
			7491: Pixel = 44;
			7492: Pixel = 48;
			7493: Pixel = 52;
			7494: Pixel = 54;
			7495: Pixel = 71;
			7496: Pixel = 109;
			7497: Pixel = 100;
			7498: Pixel = 86;
			7499: Pixel = 86;
			7500: Pixel = 62;
			7501: Pixel = 60;
			7502: Pixel = 54;
			7503: Pixel = 59;
			7504: Pixel = 61;
			7505: Pixel = 65;
			7506: Pixel = 68;
			7507: Pixel = 68;
			7508: Pixel = 66;
			7509: Pixel = 63;
			7510: Pixel = 60;
			7511: Pixel = 65;
			7512: Pixel = 63;
			7513: Pixel = 63;
			7514: Pixel = 60;
			7515: Pixel = 62;
			7516: Pixel = 59;
			7517: Pixel = 55;
			7518: Pixel = 59;
			7519: Pixel = 58;
			7520: Pixel = 60;
			7521: Pixel = 62;
			7522: Pixel = 64;
			7523: Pixel = 56;
			7524: Pixel = 58;
			7525: Pixel = 53;
			7526: Pixel = 55;
			7527: Pixel = 27;
			7528: Pixel = 135;
			7529: Pixel = 225;
			7530: Pixel = 228;
			7531: Pixel = 247;
			7532: Pixel = 245;
			7533: Pixel = 236;
			7534: Pixel = 225;
			7535: Pixel = 203;
			7536: Pixel = 220;
			7537: Pixel = 185;
			7538: Pixel = 125;
			7539: Pixel = 129;
			7540: Pixel = 130;
			7541: Pixel = 134;
			7542: Pixel = 125;
			7543: Pixel = 122;
			7544: Pixel = 114;
			7545: Pixel = 114;
			7546: Pixel = 118;
			7547: Pixel = 121;
			7548: Pixel = 127;
			7549: Pixel = 106;
			7550: Pixel = 58;
			7551: Pixel = 104;
			7552: Pixel = 110;
			7553: Pixel = 110;
			7554: Pixel = 115;
			7555: Pixel = 129;
			7556: Pixel = 145;
			7557: Pixel = 153;
			7558: Pixel = 163;
			7559: Pixel = 168;
			7560: Pixel = 180;
			7561: Pixel = 155;
			7562: Pixel = 77;
			7563: Pixel = 123;
			7564: Pixel = 154;
			7565: Pixel = 156;
			7566: Pixel = 143;
			7567: Pixel = 150;
			7568: Pixel = 209;
			7569: Pixel = 196;
			7570: Pixel = 182;
			7571: Pixel = 204;
			7572: Pixel = 227;
			7573: Pixel = 207;
			7574: Pixel = 174;
			7575: Pixel = 115;
			7576: Pixel = 99;
			7577: Pixel = 84;
			7578: Pixel = 70;
			7579: Pixel = 60;
			7580: Pixel = 52;
			7581: Pixel = 46;
			7582: Pixel = 41;
			7583: Pixel = 41;
			7584: Pixel = 39;
			7585: Pixel = 36;
			7586: Pixel = 35;
			7587: Pixel = 34;
			7588: Pixel = 37;
			7589: Pixel = 72;
			7590: Pixel = 67;
			7591: Pixel = 38;
			7592: Pixel = 41;
			7593: Pixel = 40;
			7594: Pixel = 69;
			7595: Pixel = 103;
			7596: Pixel = 126;
			7597: Pixel = 157;
			7598: Pixel = 149;
			7599: Pixel = 152;
			7600: Pixel = 62;
			7601: Pixel = 64;
			7602: Pixel = 53;
			7603: Pixel = 53;
			7604: Pixel = 56;
			7605: Pixel = 64;
			7606: Pixel = 64;
			7607: Pixel = 67;
			7608: Pixel = 67;
			7609: Pixel = 64;
			7610: Pixel = 60;
			7611: Pixel = 63;
			7612: Pixel = 63;
			7613: Pixel = 63;
			7614: Pixel = 62;
			7615: Pixel = 62;
			7616: Pixel = 60;
			7617: Pixel = 57;
			7618: Pixel = 58;
			7619: Pixel = 60;
			7620: Pixel = 61;
			7621: Pixel = 62;
			7622: Pixel = 64;
			7623: Pixel = 59;
			7624: Pixel = 60;
			7625: Pixel = 64;
			7626: Pixel = 46;
			7627: Pixel = 41;
			7628: Pixel = 88;
			7629: Pixel = 126;
			7630: Pixel = 166;
			7631: Pixel = 176;
			7632: Pixel = 202;
			7633: Pixel = 194;
			7634: Pixel = 161;
			7635: Pixel = 199;
			7636: Pixel = 222;
			7637: Pixel = 154;
			7638: Pixel = 127;
			7639: Pixel = 153;
			7640: Pixel = 136;
			7641: Pixel = 129;
			7642: Pixel = 125;
			7643: Pixel = 101;
			7644: Pixel = 86;
			7645: Pixel = 96;
			7646: Pixel = 106;
			7647: Pixel = 113;
			7648: Pixel = 117;
			7649: Pixel = 65;
			7650: Pixel = 52;
			7651: Pixel = 73;
			7652: Pixel = 86;
			7653: Pixel = 93;
			7654: Pixel = 91;
			7655: Pixel = 95;
			7656: Pixel = 107;
			7657: Pixel = 115;
			7658: Pixel = 124;
			7659: Pixel = 130;
			7660: Pixel = 133;
			7661: Pixel = 124;
			7662: Pixel = 76;
			7663: Pixel = 113;
			7664: Pixel = 141;
			7665: Pixel = 145;
			7666: Pixel = 134;
			7667: Pixel = 144;
			7668: Pixel = 169;
			7669: Pixel = 177;
			7670: Pixel = 183;
			7671: Pixel = 208;
			7672: Pixel = 238;
			7673: Pixel = 221;
			7674: Pixel = 215;
			7675: Pixel = 194;
			7676: Pixel = 198;
			7677: Pixel = 190;
			7678: Pixel = 179;
			7679: Pixel = 167;
			7680: Pixel = 151;
			7681: Pixel = 133;
			7682: Pixel = 118;
			7683: Pixel = 103;
			7684: Pixel = 86;
			7685: Pixel = 74;
			7686: Pixel = 66;
			7687: Pixel = 57;
			7688: Pixel = 54;
			7689: Pixel = 74;
			7690: Pixel = 73;
			7691: Pixel = 93;
			7692: Pixel = 102;
			7693: Pixel = 71;
			7694: Pixel = 110;
			7695: Pixel = 129;
			7696: Pixel = 129;
			7697: Pixel = 162;
			7698: Pixel = 184;
			7699: Pixel = 118;
			7700: Pixel = 58;
			7701: Pixel = 60;
			7702: Pixel = 57;
			7703: Pixel = 51;
			7704: Pixel = 51;
			7705: Pixel = 59;
			7706: Pixel = 61;
			7707: Pixel = 65;
			7708: Pixel = 64;
			7709: Pixel = 62;
			7710: Pixel = 59;
			7711: Pixel = 58;
			7712: Pixel = 61;
			7713: Pixel = 58;
			7714: Pixel = 58;
			7715: Pixel = 58;
			7716: Pixel = 60;
			7717: Pixel = 58;
			7718: Pixel = 56;
			7719: Pixel = 59;
			7720: Pixel = 60;
			7721: Pixel = 62;
			7722: Pixel = 63;
			7723: Pixel = 60;
			7724: Pixel = 62;
			7725: Pixel = 69;
			7726: Pixel = 57;
			7727: Pixel = 64;
			7728: Pixel = 62;
			7729: Pixel = 92;
			7730: Pixel = 111;
			7731: Pixel = 99;
			7732: Pixel = 101;
			7733: Pixel = 131;
			7734: Pixel = 122;
			7735: Pixel = 145;
			7736: Pixel = 171;
			7737: Pixel = 124;
			7738: Pixel = 152;
			7739: Pixel = 155;
			7740: Pixel = 135;
			7741: Pixel = 122;
			7742: Pixel = 123;
			7743: Pixel = 95;
			7744: Pixel = 66;
			7745: Pixel = 50;
			7746: Pixel = 59;
			7747: Pixel = 75;
			7748: Pixel = 64;
			7749: Pixel = 46;
			7750: Pixel = 49;
			7751: Pixel = 45;
			7752: Pixel = 55;
			7753: Pixel = 78;
			7754: Pixel = 74;
			7755: Pixel = 59;
			7756: Pixel = 67;
			7757: Pixel = 74;
			7758: Pixel = 77;
			7759: Pixel = 79;
			7760: Pixel = 88;
			7761: Pixel = 97;
			7762: Pixel = 72;
			7763: Pixel = 110;
			7764: Pixel = 118;
			7765: Pixel = 139;
			7766: Pixel = 147;
			7767: Pixel = 128;
			7768: Pixel = 130;
			7769: Pixel = 134;
			7770: Pixel = 134;
			7771: Pixel = 149;
			7772: Pixel = 182;
			7773: Pixel = 161;
			7774: Pixel = 172;
			7775: Pixel = 157;
			7776: Pixel = 172;
			7777: Pixel = 176;
			7778: Pixel = 184;
			7779: Pixel = 193;
			7780: Pixel = 199;
			7781: Pixel = 205;
			7782: Pixel = 203;
			7783: Pixel = 203;
			7784: Pixel = 189;
			7785: Pixel = 181;
			7786: Pixel = 170;
			7787: Pixel = 157;
			7788: Pixel = 151;
			7789: Pixel = 147;
			7790: Pixel = 131;
			7791: Pixel = 147;
			7792: Pixel = 195;
			7793: Pixel = 176;
			7794: Pixel = 153;
			7795: Pixel = 149;
			7796: Pixel = 169;
			7797: Pixel = 169;
			7798: Pixel = 130;
			7799: Pixel = 85;
			7800: Pixel = 54;
			7801: Pixel = 57;
			7802: Pixel = 61;
			7803: Pixel = 51;
			7804: Pixel = 50;
			7805: Pixel = 52;
			7806: Pixel = 56;
			7807: Pixel = 63;
			7808: Pixel = 64;
			7809: Pixel = 64;
			7810: Pixel = 60;
			7811: Pixel = 55;
			7812: Pixel = 61;
			7813: Pixel = 60;
			7814: Pixel = 60;
			7815: Pixel = 59;
			7816: Pixel = 63;
			7817: Pixel = 58;
			7818: Pixel = 58;
			7819: Pixel = 60;
			7820: Pixel = 60;
			7821: Pixel = 62;
			7822: Pixel = 66;
			7823: Pixel = 64;
			7824: Pixel = 65;
			7825: Pixel = 71;
			7826: Pixel = 69;
			7827: Pixel = 72;
			7828: Pixel = 67;
			7829: Pixel = 61;
			7830: Pixel = 72;
			7831: Pixel = 120;
			7832: Pixel = 166;
			7833: Pixel = 132;
			7834: Pixel = 130;
			7835: Pixel = 146;
			7836: Pixel = 132;
			7837: Pixel = 124;
			7838: Pixel = 134;
			7839: Pixel = 125;
			7840: Pixel = 125;
			7841: Pixel = 122;
			7842: Pixel = 125;
			7843: Pixel = 97;
			7844: Pixel = 69;
			7845: Pixel = 53;
			7846: Pixel = 47;
			7847: Pixel = 51;
			7848: Pixel = 49;
			7849: Pixel = 46;
			7850: Pixel = 52;
			7851: Pixel = 47;
			7852: Pixel = 47;
			7853: Pixel = 74;
			7854: Pixel = 74;
			7855: Pixel = 59;
			7856: Pixel = 65;
			7857: Pixel = 68;
			7858: Pixel = 62;
			7859: Pixel = 54;
			7860: Pixel = 54;
			7861: Pixel = 52;
			7862: Pixel = 52;
			7863: Pixel = 119;
			7864: Pixel = 151;
			7865: Pixel = 155;
			7866: Pixel = 118;
			7867: Pixel = 62;
			7868: Pixel = 73;
			7869: Pixel = 78;
			7870: Pixel = 83;
			7871: Pixel = 110;
			7872: Pixel = 123;
			7873: Pixel = 124;
			7874: Pixel = 113;
			7875: Pixel = 114;
			7876: Pixel = 125;
			7877: Pixel = 129;
			7878: Pixel = 133;
			7879: Pixel = 138;
			7880: Pixel = 144;
			7881: Pixel = 153;
			7882: Pixel = 159;
			7883: Pixel = 167;
			7884: Pixel = 173;
			7885: Pixel = 180;
			7886: Pixel = 183;
			7887: Pixel = 190;
			7888: Pixel = 198;
			7889: Pixel = 210;
			7890: Pixel = 209;
			7891: Pixel = 189;
			7892: Pixel = 211;
			7893: Pixel = 215;
			7894: Pixel = 209;
			7895: Pixel = 200;
			7896: Pixel = 232;
			7897: Pixel = 166;
			7898: Pixel = 92;
			7899: Pixel = 98;
			7900: Pixel = 52;
			7901: Pixel = 56;
			7902: Pixel = 59;
			7903: Pixel = 53;
			7904: Pixel = 47;
			7905: Pixel = 50;
			7906: Pixel = 52;
			7907: Pixel = 61;
			7908: Pixel = 66;
			7909: Pixel = 66;
			7910: Pixel = 61;
			7911: Pixel = 56;
			7912: Pixel = 61;
			7913: Pixel = 61;
			7914: Pixel = 59;
			7915: Pixel = 60;
			7916: Pixel = 62;
			7917: Pixel = 61;
			7918: Pixel = 60;
			7919: Pixel = 62;
			7920: Pixel = 61;
			7921: Pixel = 63;
			7922: Pixel = 66;
			7923: Pixel = 66;
			7924: Pixel = 66;
			7925: Pixel = 75;
			7926: Pixel = 68;
			7927: Pixel = 59;
			7928: Pixel = 77;
			7929: Pixel = 131;
			7930: Pixel = 194;
			7931: Pixel = 242;
			7932: Pixel = 232;
			7933: Pixel = 143;
			7934: Pixel = 100;
			7935: Pixel = 144;
			7936: Pixel = 129;
			7937: Pixel = 117;
			7938: Pixel = 127;
			7939: Pixel = 127;
			7940: Pixel = 126;
			7941: Pixel = 119;
			7942: Pixel = 126;
			7943: Pixel = 97;
			7944: Pixel = 74;
			7945: Pixel = 59;
			7946: Pixel = 57;
			7947: Pixel = 55;
			7948: Pixel = 55;
			7949: Pixel = 49;
			7950: Pixel = 49;
			7951: Pixel = 65;
			7952: Pixel = 52;
			7953: Pixel = 68;
			7954: Pixel = 76;
			7955: Pixel = 61;
			7956: Pixel = 67;
			7957: Pixel = 69;
			7958: Pixel = 67;
			7959: Pixel = 59;
			7960: Pixel = 55;
			7961: Pixel = 54;
			7962: Pixel = 49;
			7963: Pixel = 68;
			7964: Pixel = 92;
			7965: Pixel = 93;
			7966: Pixel = 62;
			7967: Pixel = 37;
			7968: Pixel = 38;
			7969: Pixel = 39;
			7970: Pixel = 34;
			7971: Pixel = 52;
			7972: Pixel = 73;
			7973: Pixel = 87;
			7974: Pixel = 72;
			7975: Pixel = 64;
			7976: Pixel = 67;
			7977: Pixel = 69;
			7978: Pixel = 78;
			7979: Pixel = 88;
			7980: Pixel = 91;
			7981: Pixel = 101;
			7982: Pixel = 110;
			7983: Pixel = 116;
			7984: Pixel = 123;
			7985: Pixel = 129;
			7986: Pixel = 134;
			7987: Pixel = 140;
			7988: Pixel = 145;
			7989: Pixel = 159;
			7990: Pixel = 151;
			7991: Pixel = 142;
			7992: Pixel = 169;
			7993: Pixel = 172;
			7994: Pixel = 208;
			7995: Pixel = 196;
			7996: Pixel = 192;
			7997: Pixel = 118;
			7998: Pixel = 86;
			7999: Pixel = 87;
			8000: Pixel = 51;
			8001: Pixel = 54;
			8002: Pixel = 57;
			8003: Pixel = 59;
			8004: Pixel = 50;
			8005: Pixel = 49;
			8006: Pixel = 52;
			8007: Pixel = 59;
			8008: Pixel = 64;
			8009: Pixel = 67;
			8010: Pixel = 65;
			8011: Pixel = 61;
			8012: Pixel = 58;
			8013: Pixel = 62;
			8014: Pixel = 63;
			8015: Pixel = 64;
			8016: Pixel = 65;
			8017: Pixel = 66;
			8018: Pixel = 64;
			8019: Pixel = 66;
			8020: Pixel = 66;
			8021: Pixel = 67;
			8022: Pixel = 70;
			8023: Pixel = 72;
			8024: Pixel = 65;
			8025: Pixel = 71;
			8026: Pixel = 102;
			8027: Pixel = 155;
			8028: Pixel = 219;
			8029: Pixel = 255;
			8030: Pixel = 245;
			8031: Pixel = 184;
			8032: Pixel = 128;
			8033: Pixel = 93;
			8034: Pixel = 52;
			8035: Pixel = 78;
			8036: Pixel = 135;
			8037: Pixel = 105;
			8038: Pixel = 122;
			8039: Pixel = 125;
			8040: Pixel = 120;
			8041: Pixel = 125;
			8042: Pixel = 117;
			8043: Pixel = 112;
			8044: Pixel = 102;
			8045: Pixel = 79;
			8046: Pixel = 64;
			8047: Pixel = 54;
			8048: Pixel = 55;
			8049: Pixel = 50;
			8050: Pixel = 58;
			8051: Pixel = 99;
			8052: Pixel = 66;
			8053: Pixel = 72;
			8054: Pixel = 77;
			8055: Pixel = 65;
			8056: Pixel = 68;
			8057: Pixel = 69;
			8058: Pixel = 70;
			8059: Pixel = 62;
			8060: Pixel = 56;
			8061: Pixel = 53;
			8062: Pixel = 50;
			8063: Pixel = 64;
			8064: Pixel = 79;
			8065: Pixel = 84;
			8066: Pixel = 60;
			8067: Pixel = 43;
			8068: Pixel = 42;
			8069: Pixel = 43;
			8070: Pixel = 37;
			8071: Pixel = 43;
			8072: Pixel = 44;
			8073: Pixel = 52;
			8074: Pixel = 62;
			8075: Pixel = 61;
			8076: Pixel = 55;
			8077: Pixel = 48;
			8078: Pixel = 47;
			8079: Pixel = 50;
			8080: Pixel = 53;
			8081: Pixel = 49;
			8082: Pixel = 50;
			8083: Pixel = 54;
			8084: Pixel = 59;
			8085: Pixel = 61;
			8086: Pixel = 64;
			8087: Pixel = 64;
			8088: Pixel = 75;
			8089: Pixel = 91;
			8090: Pixel = 79;
			8091: Pixel = 104;
			8092: Pixel = 110;
			8093: Pixel = 129;
			8094: Pixel = 148;
			8095: Pixel = 134;
			8096: Pixel = 100;
			8097: Pixel = 91;
			8098: Pixel = 92;
			8099: Pixel = 92;
			8100: Pixel = 56;
			8101: Pixel = 53;
			8102: Pixel = 55;
			8103: Pixel = 59;
			8104: Pixel = 51;
			8105: Pixel = 48;
			8106: Pixel = 50;
			8107: Pixel = 56;
			8108: Pixel = 64;
			8109: Pixel = 67;
			8110: Pixel = 67;
			8111: Pixel = 64;
			8112: Pixel = 61;
			8113: Pixel = 65;
			8114: Pixel = 65;
			8115: Pixel = 67;
			8116: Pixel = 66;
			8117: Pixel = 69;
			8118: Pixel = 69;
			8119: Pixel = 70;
			8120: Pixel = 73;
			8121: Pixel = 70;
			8122: Pixel = 68;
			8123: Pixel = 78;
			8124: Pixel = 119;
			8125: Pixel = 182;
			8126: Pixel = 237;
			8127: Pixel = 255;
			8128: Pixel = 246;
			8129: Pixel = 196;
			8130: Pixel = 129;
			8131: Pixel = 94;
			8132: Pixel = 92;
			8133: Pixel = 62;
			8134: Pixel = 52;
			8135: Pixel = 55;
			8136: Pixel = 121;
			8137: Pixel = 116;
			8138: Pixel = 115;
			8139: Pixel = 119;
			8140: Pixel = 126;
			8141: Pixel = 109;
			8142: Pixel = 96;
			8143: Pixel = 120;
			8144: Pixel = 127;
			8145: Pixel = 112;
			8146: Pixel = 67;
			8147: Pixel = 53;
			8148: Pixel = 48;
			8149: Pixel = 44;
			8150: Pixel = 50;
			8151: Pixel = 97;
			8152: Pixel = 96;
			8153: Pixel = 78;
			8154: Pixel = 74;
			8155: Pixel = 68;
			8156: Pixel = 72;
			8157: Pixel = 73;
			8158: Pixel = 72;
			8159: Pixel = 65;
			8160: Pixel = 57;
			8161: Pixel = 52;
			8162: Pixel = 45;
			8163: Pixel = 71;
			8164: Pixel = 108;
			8165: Pixel = 116;
			8166: Pixel = 60;
			8167: Pixel = 40;
			8168: Pixel = 41;
			8169: Pixel = 40;
			8170: Pixel = 36;
			8171: Pixel = 44;
			8172: Pixel = 48;
			8173: Pixel = 54;
			8174: Pixel = 63;
			8175: Pixel = 62;
			8176: Pixel = 60;
			8177: Pixel = 55;
			8178: Pixel = 51;
			8179: Pixel = 51;
			8180: Pixel = 55;
			8181: Pixel = 48;
			8182: Pixel = 47;
			8183: Pixel = 49;
			8184: Pixel = 47;
			8185: Pixel = 41;
			8186: Pixel = 37;
			8187: Pixel = 33;
			8188: Pixel = 45;
			8189: Pixel = 64;
			8190: Pixel = 65;
			8191: Pixel = 69;
			8192: Pixel = 85;
			8193: Pixel = 93;
			8194: Pixel = 87;
			8195: Pixel = 82;
			8196: Pixel = 74;
			8197: Pixel = 87;
			8198: Pixel = 100;
			8199: Pixel = 166;
			8200: Pixel = 63;
			8201: Pixel = 51;
			8202: Pixel = 54;
			8203: Pixel = 57;
			8204: Pixel = 59;
			8205: Pixel = 51;
			8206: Pixel = 49;
			8207: Pixel = 53;
			8208: Pixel = 63;
			8209: Pixel = 67;
			8210: Pixel = 71;
			8211: Pixel = 68;
			8212: Pixel = 64;
			8213: Pixel = 68;
			8214: Pixel = 69;
			8215: Pixel = 70;
			8216: Pixel = 69;
			8217: Pixel = 73;
			8218: Pixel = 75;
			8219: Pixel = 69;
			8220: Pixel = 68;
			8221: Pixel = 88;
			8222: Pixel = 140;
			8223: Pixel = 203;
			8224: Pixel = 249;
			8225: Pixel = 255;
			8226: Pixel = 238;
			8227: Pixel = 189;
			8228: Pixel = 128;
			8229: Pixel = 90;
			8230: Pixel = 86;
			8231: Pixel = 101;
			8232: Pixel = 77;
			8233: Pixel = 54;
			8234: Pixel = 53;
			8235: Pixel = 41;
			8236: Pixel = 68;
			8237: Pixel = 116;
			8238: Pixel = 123;
			8239: Pixel = 118;
			8240: Pixel = 112;
			8241: Pixel = 64;
			8242: Pixel = 97;
			8243: Pixel = 162;
			8244: Pixel = 91;
			8245: Pixel = 90;
			8246: Pixel = 68;
			8247: Pixel = 52;
			8248: Pixel = 45;
			8249: Pixel = 48;
			8250: Pixel = 38;
			8251: Pixel = 82;
			8252: Pixel = 93;
			8253: Pixel = 64;
			8254: Pixel = 72;
			8255: Pixel = 74;
			8256: Pixel = 77;
			8257: Pixel = 79;
			8258: Pixel = 79;
			8259: Pixel = 74;
			8260: Pixel = 59;
			8261: Pixel = 52;
			8262: Pixel = 45;
			8263: Pixel = 72;
			8264: Pixel = 133;
			8265: Pixel = 138;
			8266: Pixel = 61;
			8267: Pixel = 38;
			8268: Pixel = 42;
			8269: Pixel = 40;
			8270: Pixel = 34;
			8271: Pixel = 43;
			8272: Pixel = 45;
			8273: Pixel = 52;
			8274: Pixel = 58;
			8275: Pixel = 60;
			8276: Pixel = 61;
			8277: Pixel = 62;
			8278: Pixel = 53;
			8279: Pixel = 52;
			8280: Pixel = 53;
			8281: Pixel = 48;
			8282: Pixel = 47;
			8283: Pixel = 48;
			8284: Pixel = 46;
			8285: Pixel = 43;
			8286: Pixel = 41;
			8287: Pixel = 36;
			8288: Pixel = 49;
			8289: Pixel = 64;
			8290: Pixel = 70;
			8291: Pixel = 38;
			8292: Pixel = 52;
			8293: Pixel = 79;
			8294: Pixel = 95;
			8295: Pixel = 95;
			8296: Pixel = 56;
			8297: Pixel = 69;
			8298: Pixel = 116;
			8299: Pixel = 152;
			8300: Pixel = 62;
			8301: Pixel = 53;
			8302: Pixel = 54;
			8303: Pixel = 59;
			8304: Pixel = 62;
			8305: Pixel = 51;
			8306: Pixel = 46;
			8307: Pixel = 54;
			8308: Pixel = 60;
			8309: Pixel = 70;
			8310: Pixel = 71;
			8311: Pixel = 72;
			8312: Pixel = 69;
			8313: Pixel = 71;
			8314: Pixel = 75;
			8315: Pixel = 77;
			8316: Pixel = 78;
			8317: Pixel = 74;
			8318: Pixel = 74;
			8319: Pixel = 100;
			8320: Pixel = 160;
			8321: Pixel = 222;
			8322: Pixel = 255;
			8323: Pixel = 255;
			8324: Pixel = 227;
			8325: Pixel = 178;
			8326: Pixel = 126;
			8327: Pixel = 86;
			8328: Pixel = 69;
			8329: Pixel = 92;
			8330: Pixel = 112;
			8331: Pixel = 87;
			8332: Pixel = 63;
			8333: Pixel = 58;
			8334: Pixel = 46;
			8335: Pixel = 40;
			8336: Pixel = 36;
			8337: Pixel = 51;
			8338: Pixel = 67;
			8339: Pixel = 61;
			8340: Pixel = 77;
			8341: Pixel = 70;
			8342: Pixel = 117;
			8343: Pixel = 186;
			8344: Pixel = 88;
			8345: Pixel = 71;
			8346: Pixel = 67;
			8347: Pixel = 48;
			8348: Pixel = 45;
			8349: Pixel = 49;
			8350: Pixel = 43;
			8351: Pixel = 48;
			8352: Pixel = 59;
			8353: Pixel = 57;
			8354: Pixel = 70;
			8355: Pixel = 79;
			8356: Pixel = 81;
			8357: Pixel = 81;
			8358: Pixel = 82;
			8359: Pixel = 77;
			8360: Pixel = 63;
			8361: Pixel = 52;
			8362: Pixel = 44;
			8363: Pixel = 70;
			8364: Pixel = 124;
			8365: Pixel = 127;
			8366: Pixel = 60;
			8367: Pixel = 39;
			8368: Pixel = 42;
			8369: Pixel = 37;
			8370: Pixel = 31;
			8371: Pixel = 42;
			8372: Pixel = 43;
			8373: Pixel = 49;
			8374: Pixel = 56;
			8375: Pixel = 58;
			8376: Pixel = 60;
			8377: Pixel = 66;
			8378: Pixel = 57;
			8379: Pixel = 49;
			8380: Pixel = 48;
			8381: Pixel = 45;
			8382: Pixel = 45;
			8383: Pixel = 47;
			8384: Pixel = 45;
			8385: Pixel = 43;
			8386: Pixel = 39;
			8387: Pixel = 35;
			8388: Pixel = 52;
			8389: Pixel = 65;
			8390: Pixel = 68;
			8391: Pixel = 38;
			8392: Pixel = 36;
			8393: Pixel = 97;
			8394: Pixel = 139;
			8395: Pixel = 81;
			8396: Pixel = 47;
			8397: Pixel = 64;
			8398: Pixel = 94;
			8399: Pixel = 145;
			8400: Pixel = 62;
			8401: Pixel = 58;
			8402: Pixel = 55;
			8403: Pixel = 63;
			8404: Pixel = 62;
			8405: Pixel = 59;
			8406: Pixel = 52;
			8407: Pixel = 54;
			8408: Pixel = 60;
			8409: Pixel = 70;
			8410: Pixel = 74;
			8411: Pixel = 78;
			8412: Pixel = 76;
			8413: Pixel = 76;
			8414: Pixel = 79;
			8415: Pixel = 75;
			8416: Pixel = 80;
			8417: Pixel = 120;
			8418: Pixel = 183;
			8419: Pixel = 236;
			8420: Pixel = 255;
			8421: Pixel = 250;
			8422: Pixel = 211;
			8423: Pixel = 158;
			8424: Pixel = 108;
			8425: Pixel = 79;
			8426: Pixel = 79;
			8427: Pixel = 95;
			8428: Pixel = 120;
			8429: Pixel = 120;
			8430: Pixel = 86;
			8431: Pixel = 74;
			8432: Pixel = 67;
			8433: Pixel = 53;
			8434: Pixel = 41;
			8435: Pixel = 40;
			8436: Pixel = 37;
			8437: Pixel = 42;
			8438: Pixel = 40;
			8439: Pixel = 44;
			8440: Pixel = 55;
			8441: Pixel = 63;
			8442: Pixel = 109;
			8443: Pixel = 124;
			8444: Pixel = 88;
			8445: Pixel = 77;
			8446: Pixel = 68;
			8447: Pixel = 50;
			8448: Pixel = 47;
			8449: Pixel = 51;
			8450: Pixel = 48;
			8451: Pixel = 45;
			8452: Pixel = 57;
			8453: Pixel = 72;
			8454: Pixel = 72;
			8455: Pixel = 81;
			8456: Pixel = 84;
			8457: Pixel = 84;
			8458: Pixel = 81;
			8459: Pixel = 77;
			8460: Pixel = 68;
			8461: Pixel = 52;
			8462: Pixel = 45;
			8463: Pixel = 72;
			8464: Pixel = 119;
			8465: Pixel = 127;
			8466: Pixel = 61;
			8467: Pixel = 39;
			8468: Pixel = 44;
			8469: Pixel = 39;
			8470: Pixel = 33;
			8471: Pixel = 42;
			8472: Pixel = 45;
			8473: Pixel = 48;
			8474: Pixel = 55;
			8475: Pixel = 59;
			8476: Pixel = 59;
			8477: Pixel = 64;
			8478: Pixel = 61;
			8479: Pixel = 54;
			8480: Pixel = 47;
			8481: Pixel = 50;
			8482: Pixel = 63;
			8483: Pixel = 47;
			8484: Pixel = 45;
			8485: Pixel = 40;
			8486: Pixel = 38;
			8487: Pixel = 38;
			8488: Pixel = 52;
			8489: Pixel = 67;
			8490: Pixel = 69;
			8491: Pixel = 43;
			8492: Pixel = 39;
			8493: Pixel = 64;
			8494: Pixel = 106;
			8495: Pixel = 66;
			8496: Pixel = 53;
			8497: Pixel = 59;
			8498: Pixel = 95;
			8499: Pixel = 128;
			8500: Pixel = 59;
			8501: Pixel = 61;
			8502: Pixel = 56;
			8503: Pixel = 63;
			8504: Pixel = 61;
			8505: Pixel = 65;
			8506: Pixel = 57;
			8507: Pixel = 56;
			8508: Pixel = 60;
			8509: Pixel = 71;
			8510: Pixel = 80;
			8511: Pixel = 84;
			8512: Pixel = 79;
			8513: Pixel = 70;
			8514: Pixel = 87;
			8515: Pixel = 132;
			8516: Pixel = 194;
			8517: Pixel = 244;
			8518: Pixel = 255;
			8519: Pixel = 245;
			8520: Pixel = 198;
			8521: Pixel = 140;
			8522: Pixel = 95;
			8523: Pixel = 75;
			8524: Pixel = 72;
			8525: Pixel = 83;
			8526: Pixel = 123;
			8527: Pixel = 112;
			8528: Pixel = 100;
			8529: Pixel = 76;
			8530: Pixel = 74;
			8531: Pixel = 79;
			8532: Pixel = 57;
			8533: Pixel = 38;
			8534: Pixel = 40;
			8535: Pixel = 39;
			8536: Pixel = 35;
			8537: Pixel = 36;
			8538: Pixel = 35;
			8539: Pixel = 41;
			8540: Pixel = 48;
			8541: Pixel = 60;
			8542: Pixel = 67;
			8543: Pixel = 110;
			8544: Pixel = 95;
			8545: Pixel = 91;
			8546: Pixel = 76;
			8547: Pixel = 54;
			8548: Pixel = 52;
			8549: Pixel = 51;
			8550: Pixel = 50;
			8551: Pixel = 50;
			8552: Pixel = 65;
			8553: Pixel = 72;
			8554: Pixel = 76;
			8555: Pixel = 81;
			8556: Pixel = 82;
			8557: Pixel = 82;
			8558: Pixel = 79;
			8559: Pixel = 80;
			8560: Pixel = 79;
			8561: Pixel = 57;
			8562: Pixel = 44;
			8563: Pixel = 71;
			8564: Pixel = 118;
			8565: Pixel = 125;
			8566: Pixel = 60;
			8567: Pixel = 40;
			8568: Pixel = 45;
			8569: Pixel = 38;
			8570: Pixel = 32;
			8571: Pixel = 41;
			8572: Pixel = 44;
			8573: Pixel = 48;
			8574: Pixel = 54;
			8575: Pixel = 58;
			8576: Pixel = 59;
			8577: Pixel = 60;
			8578: Pixel = 58;
			8579: Pixel = 55;
			8580: Pixel = 46;
			8581: Pixel = 49;
			8582: Pixel = 64;
			8583: Pixel = 44;
			8584: Pixel = 42;
			8585: Pixel = 39;
			8586: Pixel = 37;
			8587: Pixel = 39;
			8588: Pixel = 47;
			8589: Pixel = 63;
			8590: Pixel = 71;
			8591: Pixel = 45;
			8592: Pixel = 44;
			8593: Pixel = 49;
			8594: Pixel = 52;
			8595: Pixel = 60;
			8596: Pixel = 57;
			8597: Pixel = 59;
			8598: Pixel = 100;
			8599: Pixel = 117;
			8600: Pixel = 58;
			8601: Pixel = 63;
			8602: Pixel = 59;
			8603: Pixel = 63;
			8604: Pixel = 65;
			8605: Pixel = 67;
			8606: Pixel = 64;
			8607: Pixel = 60;
			8608: Pixel = 65;
			8609: Pixel = 78;
			8610: Pixel = 79;
			8611: Pixel = 78;
			8612: Pixel = 99;
			8613: Pixel = 149;
			8614: Pixel = 208;
			8615: Pixel = 251;
			8616: Pixel = 255;
			8617: Pixel = 241;
			8618: Pixel = 195;
			8619: Pixel = 133;
			8620: Pixel = 88;
			8621: Pixel = 73;
			8622: Pixel = 74;
			8623: Pixel = 74;
			8624: Pixel = 69;
			8625: Pixel = 78;
			8626: Pixel = 95;
			8627: Pixel = 73;
			8628: Pixel = 67;
			8629: Pixel = 71;
			8630: Pixel = 73;
			8631: Pixel = 60;
			8632: Pixel = 38;
			8633: Pixel = 37;
			8634: Pixel = 38;
			8635: Pixel = 36;
			8636: Pixel = 36;
			8637: Pixel = 33;
			8638: Pixel = 34;
			8639: Pixel = 40;
			8640: Pixel = 48;
			8641: Pixel = 56;
			8642: Pixel = 63;
			8643: Pixel = 107;
			8644: Pixel = 107;
			8645: Pixel = 102;
			8646: Pixel = 86;
			8647: Pixel = 64;
			8648: Pixel = 53;
			8649: Pixel = 49;
			8650: Pixel = 53;
			8651: Pixel = 56;
			8652: Pixel = 65;
			8653: Pixel = 72;
			8654: Pixel = 78;
			8655: Pixel = 82;
			8656: Pixel = 84;
			8657: Pixel = 84;
			8658: Pixel = 81;
			8659: Pixel = 80;
			8660: Pixel = 85;
			8661: Pixel = 71;
			8662: Pixel = 47;
			8663: Pixel = 71;
			8664: Pixel = 115;
			8665: Pixel = 124;
			8666: Pixel = 61;
			8667: Pixel = 40;
			8668: Pixel = 45;
			8669: Pixel = 36;
			8670: Pixel = 33;
			8671: Pixel = 41;
			8672: Pixel = 44;
			8673: Pixel = 48;
			8674: Pixel = 53;
			8675: Pixel = 56;
			8676: Pixel = 56;
			8677: Pixel = 57;
			8678: Pixel = 57;
			8679: Pixel = 54;
			8680: Pixel = 49;
			8681: Pixel = 46;
			8682: Pixel = 42;
			8683: Pixel = 40;
			8684: Pixel = 38;
			8685: Pixel = 38;
			8686: Pixel = 39;
			8687: Pixel = 37;
			8688: Pixel = 47;
			8689: Pixel = 59;
			8690: Pixel = 75;
			8691: Pixel = 53;
			8692: Pixel = 48;
			8693: Pixel = 53;
			8694: Pixel = 54;
			8695: Pixel = 62;
			8696: Pixel = 63;
			8697: Pixel = 76;
			8698: Pixel = 120;
			8699: Pixel = 145;
			8700: Pixel = 62;
			8701: Pixel = 61;
			8702: Pixel = 65;
			8703: Pixel = 58;
			8704: Pixel = 68;
			8705: Pixel = 67;
			8706: Pixel = 69;
			8707: Pixel = 66;
			8708: Pixel = 71;
			8709: Pixel = 80;
			8710: Pixel = 111;
			8711: Pixel = 164;
			8712: Pixel = 223;
			8713: Pixel = 255;
			8714: Pixel = 255;
			8715: Pixel = 236;
			8716: Pixel = 190;
			8717: Pixel = 129;
			8718: Pixel = 85;
			8719: Pixel = 74;
			8720: Pixel = 71;
			8721: Pixel = 74;
			8722: Pixel = 73;
			8723: Pixel = 71;
			8724: Pixel = 67;
			8725: Pixel = 66;
			8726: Pixel = 65;
			8727: Pixel = 68;
			8728: Pixel = 66;
			8729: Pixel = 60;
			8730: Pixel = 64;
			8731: Pixel = 42;
			8732: Pixel = 32;
			8733: Pixel = 42;
			8734: Pixel = 44;
			8735: Pixel = 34;
			8736: Pixel = 34;
			8737: Pixel = 30;
			8738: Pixel = 30;
			8739: Pixel = 33;
			8740: Pixel = 44;
			8741: Pixel = 51;
			8742: Pixel = 65;
			8743: Pixel = 103;
			8744: Pixel = 108;
			8745: Pixel = 110;
			8746: Pixel = 96;
			8747: Pixel = 73;
			8748: Pixel = 51;
			8749: Pixel = 49;
			8750: Pixel = 50;
			8751: Pixel = 58;
			8752: Pixel = 68;
			8753: Pixel = 73;
			8754: Pixel = 78;
			8755: Pixel = 84;
			8756: Pixel = 84;
			8757: Pixel = 85;
			8758: Pixel = 82;
			8759: Pixel = 79;
			8760: Pixel = 81;
			8761: Pixel = 80;
			8762: Pixel = 50;
			8763: Pixel = 71;
			8764: Pixel = 112;
			8765: Pixel = 126;
			8766: Pixel = 60;
			8767: Pixel = 40;
			8768: Pixel = 46;
			8769: Pixel = 39;
			8770: Pixel = 33;
			8771: Pixel = 38;
			8772: Pixel = 44;
			8773: Pixel = 48;
			8774: Pixel = 51;
			8775: Pixel = 53;
			8776: Pixel = 55;
			8777: Pixel = 52;
			8778: Pixel = 55;
			8779: Pixel = 51;
			8780: Pixel = 42;
			8781: Pixel = 36;
			8782: Pixel = 37;
			8783: Pixel = 43;
			8784: Pixel = 37;
			8785: Pixel = 37;
			8786: Pixel = 39;
			8787: Pixel = 34;
			8788: Pixel = 44;
			8789: Pixel = 60;
			8790: Pixel = 75;
			8791: Pixel = 65;
			8792: Pixel = 47;
			8793: Pixel = 55;
			8794: Pixel = 57;
			8795: Pixel = 62;
			8796: Pixel = 67;
			8797: Pixel = 69;
			8798: Pixel = 97;
			8799: Pixel = 128;
			8800: Pixel = 69;
			8801: Pixel = 63;
			8802: Pixel = 70;
			8803: Pixel = 63;
			8804: Pixel = 73;
			8805: Pixel = 72;
			8806: Pixel = 66;
			8807: Pixel = 67;
			8808: Pixel = 107;
			8809: Pixel = 185;
			8810: Pixel = 236;
			8811: Pixel = 255;
			8812: Pixel = 255;
			8813: Pixel = 228;
			8814: Pixel = 179;
			8815: Pixel = 123;
			8816: Pixel = 87;
			8817: Pixel = 75;
			8818: Pixel = 77;
			8819: Pixel = 78;
			8820: Pixel = 71;
			8821: Pixel = 69;
			8822: Pixel = 68;
			8823: Pixel = 69;
			8824: Pixel = 65;
			8825: Pixel = 65;
			8826: Pixel = 66;
			8827: Pixel = 57;
			8828: Pixel = 44;
			8829: Pixel = 32;
			8830: Pixel = 51;
			8831: Pixel = 49;
			8832: Pixel = 31;
			8833: Pixel = 35;
			8834: Pixel = 45;
			8835: Pixel = 37;
			8836: Pixel = 36;
			8837: Pixel = 36;
			8838: Pixel = 27;
			8839: Pixel = 30;
			8840: Pixel = 41;
			8841: Pixel = 52;
			8842: Pixel = 68;
			8843: Pixel = 98;
			8844: Pixel = 109;
			8845: Pixel = 116;
			8846: Pixel = 108;
			8847: Pixel = 86;
			8848: Pixel = 60;
			8849: Pixel = 47;
			8850: Pixel = 50;
			8851: Pixel = 65;
			8852: Pixel = 72;
			8853: Pixel = 73;
			8854: Pixel = 82;
			8855: Pixel = 85;
			8856: Pixel = 84;
			8857: Pixel = 85;
			8858: Pixel = 86;
			8859: Pixel = 87;
			8860: Pixel = 82;
			8861: Pixel = 82;
			8862: Pixel = 58;
			8863: Pixel = 71;
			8864: Pixel = 111;
			8865: Pixel = 125;
			8866: Pixel = 62;
			8867: Pixel = 42;
			8868: Pixel = 46;
			8869: Pixel = 41;
			8870: Pixel = 34;
			8871: Pixel = 39;
			8872: Pixel = 45;
			8873: Pixel = 52;
			8874: Pixel = 51;
			8875: Pixel = 52;
			8876: Pixel = 54;
			8877: Pixel = 56;
			8878: Pixel = 50;
			8879: Pixel = 40;
			8880: Pixel = 34;
			8881: Pixel = 36;
			8882: Pixel = 49;
			8883: Pixel = 53;
			8884: Pixel = 39;
			8885: Pixel = 38;
			8886: Pixel = 39;
			8887: Pixel = 38;
			8888: Pixel = 45;
			8889: Pixel = 63;
			8890: Pixel = 69;
			8891: Pixel = 84;
			8892: Pixel = 51;
			8893: Pixel = 57;
			8894: Pixel = 59;
			8895: Pixel = 65;
			8896: Pixel = 70;
			8897: Pixel = 72;
			8898: Pixel = 69;
			8899: Pixel = 71;
			8900: Pixel = 75;
			8901: Pixel = 67;
			8902: Pixel = 72;
			8903: Pixel = 66;
			8904: Pixel = 62;
			8905: Pixel = 69;
			8906: Pixel = 103;
			8907: Pixel = 166;
			8908: Pixel = 233;
			8909: Pixel = 255;
			8910: Pixel = 247;
			8911: Pixel = 218;
			8912: Pixel = 168;
			8913: Pixel = 115;
			8914: Pixel = 81;
			8915: Pixel = 79;
			8916: Pixel = 80;
			8917: Pixel = 76;
			8918: Pixel = 74;
			8919: Pixel = 73;
			8920: Pixel = 67;
			8921: Pixel = 64;
			8922: Pixel = 67;
			8923: Pixel = 66;
			8924: Pixel = 61;
			8925: Pixel = 61;
			8926: Pixel = 51;
			8927: Pixel = 31;
			8928: Pixel = 28;
			8929: Pixel = 24;
			8930: Pixel = 42;
			8931: Pixel = 55;
			8932: Pixel = 27;
			8933: Pixel = 37;
			8934: Pixel = 60;
			8935: Pixel = 41;
			8936: Pixel = 37;
			8937: Pixel = 42;
			8938: Pixel = 34;
			8939: Pixel = 29;
			8940: Pixel = 38;
			8941: Pixel = 55;
			8942: Pixel = 71;
			8943: Pixel = 96;
			8944: Pixel = 110;
			8945: Pixel = 120;
			8946: Pixel = 119;
			8947: Pixel = 98;
			8948: Pixel = 71;
			8949: Pixel = 46;
			8950: Pixel = 51;
			8951: Pixel = 65;
			8952: Pixel = 75;
			8953: Pixel = 74;
			8954: Pixel = 84;
			8955: Pixel = 86;
			8956: Pixel = 87;
			8957: Pixel = 85;
			8958: Pixel = 86;
			8959: Pixel = 88;
			8960: Pixel = 87;
			8961: Pixel = 88;
			8962: Pixel = 71;
			8963: Pixel = 73;
			8964: Pixel = 111;
			8965: Pixel = 122;
			8966: Pixel = 61;
			8967: Pixel = 43;
			8968: Pixel = 47;
			8969: Pixel = 39;
			8970: Pixel = 36;
			8971: Pixel = 40;
			8972: Pixel = 47;
			8973: Pixel = 56;
			8974: Pixel = 54;
			8975: Pixel = 49;
			8976: Pixel = 51;
			8977: Pixel = 44;
			8978: Pixel = 38;
			8979: Pixel = 38;
			8980: Pixel = 41;
			8981: Pixel = 42;
			8982: Pixel = 64;
			8983: Pixel = 62;
			8984: Pixel = 38;
			8985: Pixel = 40;
			8986: Pixel = 40;
			8987: Pixel = 39;
			8988: Pixel = 39;
			8989: Pixel = 61;
			8990: Pixel = 58;
			8991: Pixel = 99;
			8992: Pixel = 57;
			8993: Pixel = 61;
			8994: Pixel = 63;
			8995: Pixel = 68;
			8996: Pixel = 71;
			8997: Pixel = 74;
			8998: Pixel = 76;
			8999: Pixel = 77;
			9000: Pixel = 82;
			9001: Pixel = 66;
			9002: Pixel = 63;
			9003: Pixel = 84;
			9004: Pixel = 128;
			9005: Pixel = 192;
			9006: Pixel = 241;
			9007: Pixel = 254;
			9008: Pixel = 231;
			9009: Pixel = 195;
			9010: Pixel = 150;
			9011: Pixel = 97;
			9012: Pixel = 76;
			9013: Pixel = 79;
			9014: Pixel = 74;
			9015: Pixel = 77;
			9016: Pixel = 77;
			9017: Pixel = 73;
			9018: Pixel = 72;
			9019: Pixel = 69;
			9020: Pixel = 63;
			9021: Pixel = 59;
			9022: Pixel = 63;
			9023: Pixel = 61;
			9024: Pixel = 58;
			9025: Pixel = 59;
			9026: Pixel = 46;
			9027: Pixel = 24;
			9028: Pixel = 28;
			9029: Pixel = 23;
			9030: Pixel = 35;
			9031: Pixel = 52;
			9032: Pixel = 28;
			9033: Pixel = 45;
			9034: Pixel = 57;
			9035: Pixel = 41;
			9036: Pixel = 39;
			9037: Pixel = 41;
			9038: Pixel = 41;
			9039: Pixel = 31;
			9040: Pixel = 36;
			9041: Pixel = 55;
			9042: Pixel = 76;
			9043: Pixel = 96;
			9044: Pixel = 105;
			9045: Pixel = 116;
			9046: Pixel = 126;
			9047: Pixel = 105;
			9048: Pixel = 81;
			9049: Pixel = 51;
			9050: Pixel = 45;
			9051: Pixel = 65;
			9052: Pixel = 79;
			9053: Pixel = 77;
			9054: Pixel = 84;
			9055: Pixel = 86;
			9056: Pixel = 87;
			9057: Pixel = 88;
			9058: Pixel = 89;
			9059: Pixel = 86;
			9060: Pixel = 86;
			9061: Pixel = 87;
			9062: Pixel = 80;
			9063: Pixel = 79;
			9064: Pixel = 110;
			9065: Pixel = 121;
			9066: Pixel = 64;
			9067: Pixel = 46;
			9068: Pixel = 46;
			9069: Pixel = 40;
			9070: Pixel = 38;
			9071: Pixel = 42;
			9072: Pixel = 53;
			9073: Pixel = 57;
			9074: Pixel = 50;
			9075: Pixel = 40;
			9076: Pixel = 39;
			9077: Pixel = 43;
			9078: Pixel = 50;
			9079: Pixel = 51;
			9080: Pixel = 52;
			9081: Pixel = 49;
			9082: Pixel = 56;
			9083: Pixel = 56;
			9084: Pixel = 38;
			9085: Pixel = 43;
			9086: Pixel = 39;
			9087: Pixel = 38;
			9088: Pixel = 37;
			9089: Pixel = 60;
			9090: Pixel = 50;
			9091: Pixel = 99;
			9092: Pixel = 79;
			9093: Pixel = 58;
			9094: Pixel = 66;
			9095: Pixel = 71;
			9096: Pixel = 73;
			9097: Pixel = 75;
			9098: Pixel = 77;
			9099: Pixel = 78;
			9100: Pixel = 87;
			9101: Pixel = 112;
			9102: Pixel = 165;
			9103: Pixel = 223;
			9104: Pixel = 254;
			9105: Pixel = 248;
			9106: Pixel = 215;
			9107: Pixel = 172;
			9108: Pixel = 149;
			9109: Pixel = 143;
			9110: Pixel = 89;
			9111: Pixel = 63;
			9112: Pixel = 72;
			9113: Pixel = 75;
			9114: Pixel = 69;
			9115: Pixel = 68;
			9116: Pixel = 71;
			9117: Pixel = 66;
			9118: Pixel = 65;
			9119: Pixel = 65;
			9120: Pixel = 62;
			9121: Pixel = 56;
			9122: Pixel = 58;
			9123: Pixel = 57;
			9124: Pixel = 55;
			9125: Pixel = 56;
			9126: Pixel = 47;
			9127: Pixel = 23;
			9128: Pixel = 23;
			9129: Pixel = 22;
			9130: Pixel = 25;
			9131: Pixel = 44;
			9132: Pixel = 31;
			9133: Pixel = 40;
			9134: Pixel = 44;
			9135: Pixel = 39;
			9136: Pixel = 39;
			9137: Pixel = 36;
			9138: Pixel = 34;
			9139: Pixel = 27;
			9140: Pixel = 33;
			9141: Pixel = 54;
			9142: Pixel = 77;
			9143: Pixel = 95;
			9144: Pixel = 102;
			9145: Pixel = 111;
			9146: Pixel = 130;
			9147: Pixel = 114;
			9148: Pixel = 89;
			9149: Pixel = 60;
			9150: Pixel = 44;
			9151: Pixel = 64;
			9152: Pixel = 78;
			9153: Pixel = 79;
			9154: Pixel = 78;
			9155: Pixel = 86;
			9156: Pixel = 89;
			9157: Pixel = 88;
			9158: Pixel = 91;
			9159: Pixel = 89;
			9160: Pixel = 87;
			9161: Pixel = 86;
			9162: Pixel = 85;
			9163: Pixel = 82;
			9164: Pixel = 107;
			9165: Pixel = 120;
			9166: Pixel = 64;
			9167: Pixel = 49;
			9168: Pixel = 46;
			9169: Pixel = 45;
			9170: Pixel = 39;
			9171: Pixel = 42;
			9172: Pixel = 45;
			9173: Pixel = 42;
			9174: Pixel = 38;
			9175: Pixel = 41;
			9176: Pixel = 43;
			9177: Pixel = 51;
			9178: Pixel = 56;
			9179: Pixel = 60;
			9180: Pixel = 58;
			9181: Pixel = 55;
			9182: Pixel = 55;
			9183: Pixel = 46;
			9184: Pixel = 39;
			9185: Pixel = 47;
			9186: Pixel = 42;
			9187: Pixel = 42;
			9188: Pixel = 41;
			9189: Pixel = 61;
			9190: Pixel = 64;
			9191: Pixel = 78;
			9192: Pixel = 112;
			9193: Pixel = 56;
			9194: Pixel = 67;
			9195: Pixel = 74;
			9196: Pixel = 75;
			9197: Pixel = 76;
			9198: Pixel = 82;
			9199: Pixel = 119;
			9200: Pixel = 200;
			9201: Pixel = 246;
			9202: Pixel = 255;
			9203: Pixel = 238;
			9204: Pixel = 192;
			9205: Pixel = 151;
			9206: Pixel = 123;
			9207: Pixel = 115;
			9208: Pixel = 112;
			9209: Pixel = 111;
			9210: Pixel = 79;
			9211: Pixel = 64;
			9212: Pixel = 63;
			9213: Pixel = 67;
			9214: Pixel = 66;
			9215: Pixel = 61;
			9216: Pixel = 68;
			9217: Pixel = 67;
			9218: Pixel = 64;
			9219: Pixel = 62;
			9220: Pixel = 61;
			9221: Pixel = 55;
			9222: Pixel = 56;
			9223: Pixel = 56;
			9224: Pixel = 54;
			9225: Pixel = 52;
			9226: Pixel = 52;
			9227: Pixel = 28;
			9228: Pixel = 24;
			9229: Pixel = 23;
			9230: Pixel = 22;
			9231: Pixel = 49;
			9232: Pixel = 31;
			9233: Pixel = 38;
			9234: Pixel = 44;
			9235: Pixel = 40;
			9236: Pixel = 41;
			9237: Pixel = 34;
			9238: Pixel = 34;
			9239: Pixel = 34;
			9240: Pixel = 31;
			9241: Pixel = 56;
			9242: Pixel = 77;
			9243: Pixel = 94;
			9244: Pixel = 104;
			9245: Pixel = 107;
			9246: Pixel = 128;
			9247: Pixel = 125;
			9248: Pixel = 99;
			9249: Pixel = 72;
			9250: Pixel = 46;
			9251: Pixel = 61;
			9252: Pixel = 80;
			9253: Pixel = 80;
			9254: Pixel = 74;
			9255: Pixel = 85;
			9256: Pixel = 90;
			9257: Pixel = 90;
			9258: Pixel = 90;
			9259: Pixel = 86;
			9260: Pixel = 90;
			9261: Pixel = 84;
			9262: Pixel = 82;
			9263: Pixel = 87;
			9264: Pixel = 108;
			9265: Pixel = 116;
			9266: Pixel = 62;
			9267: Pixel = 48;
			9268: Pixel = 48;
			9269: Pixel = 44;
			9270: Pixel = 39;
			9271: Pixel = 43;
			9272: Pixel = 46;
			9273: Pixel = 39;
			9274: Pixel = 42;
			9275: Pixel = 49;
			9276: Pixel = 47;
			9277: Pixel = 56;
			9278: Pixel = 67;
			9279: Pixel = 60;
			9280: Pixel = 58;
			9281: Pixel = 63;
			9282: Pixel = 76;
			9283: Pixel = 66;
			9284: Pixel = 46;
			9285: Pixel = 50;
			9286: Pixel = 46;
			9287: Pixel = 44;
			9288: Pixel = 44;
			9289: Pixel = 64;
			9290: Pixel = 83;
			9291: Pixel = 57;
			9292: Pixel = 122;
			9293: Pixel = 74;
			9294: Pixel = 68;
			9295: Pixel = 81;
			9296: Pixel = 78;
			9297: Pixel = 89;
			9298: Pixel = 145;
			9299: Pixel = 218;
			9300: Pixel = 252;
			9301: Pixel = 224;
			9302: Pixel = 178;
			9303: Pixel = 129;
			9304: Pixel = 113;
			9305: Pixel = 102;
			9306: Pixel = 96;
			9307: Pixel = 91;
			9308: Pixel = 93;
			9309: Pixel = 96;
			9310: Pixel = 65;
			9311: Pixel = 64;
			9312: Pixel = 57;
			9313: Pixel = 62;
			9314: Pixel = 62;
			9315: Pixel = 57;
			9316: Pixel = 63;
			9317: Pixel = 63;
			9318: Pixel = 61;
			9319: Pixel = 61;
			9320: Pixel = 57;
			9321: Pixel = 56;
			9322: Pixel = 55;
			9323: Pixel = 55;
			9324: Pixel = 52;
			9325: Pixel = 52;
			9326: Pixel = 54;
			9327: Pixel = 30;
			9328: Pixel = 21;
			9329: Pixel = 22;
			9330: Pixel = 19;
			9331: Pixel = 44;
			9332: Pixel = 36;
			9333: Pixel = 22;
			9334: Pixel = 40;
			9335: Pixel = 40;
			9336: Pixel = 41;
			9337: Pixel = 34;
			9338: Pixel = 36;
			9339: Pixel = 38;
			9340: Pixel = 28;
			9341: Pixel = 51;
			9342: Pixel = 74;
			9343: Pixel = 93;
			9344: Pixel = 107;
			9345: Pixel = 102;
			9346: Pixel = 124;
			9347: Pixel = 130;
			9348: Pixel = 107;
			9349: Pixel = 83;
			9350: Pixel = 51;
			9351: Pixel = 52;
			9352: Pixel = 77;
			9353: Pixel = 79;
			9354: Pixel = 72;
			9355: Pixel = 78;
			9356: Pixel = 82;
			9357: Pixel = 86;
			9358: Pixel = 84;
			9359: Pixel = 85;
			9360: Pixel = 85;
			9361: Pixel = 83;
			9362: Pixel = 75;
			9363: Pixel = 84;
			9364: Pixel = 108;
			9365: Pixel = 116;
			9366: Pixel = 65;
			9367: Pixel = 42;
			9368: Pixel = 39;
			9369: Pixel = 39;
			9370: Pixel = 39;
			9371: Pixel = 44;
			9372: Pixel = 56;
			9373: Pixel = 45;
			9374: Pixel = 42;
			9375: Pixel = 47;
			9376: Pixel = 49;
			9377: Pixel = 60;
			9378: Pixel = 64;
			9379: Pixel = 66;
			9380: Pixel = 76;
			9381: Pixel = 75;
			9382: Pixel = 80;
			9383: Pixel = 69;
			9384: Pixel = 63;
			9385: Pixel = 49;
			9386: Pixel = 45;
			9387: Pixel = 45;
			9388: Pixel = 47;
			9389: Pixel = 62;
			9390: Pixel = 86;
			9391: Pixel = 66;
			9392: Pixel = 102;
			9393: Pixel = 116;
			9394: Pixel = 65;
			9395: Pixel = 85;
			9396: Pixel = 113;
			9397: Pixel = 172;
			9398: Pixel = 232;
			9399: Pixel = 249;
			9400: Pixel = 168;
			9401: Pixel = 136;
			9402: Pixel = 93;
			9403: Pixel = 73;
			9404: Pixel = 96;
			9405: Pixel = 90;
			9406: Pixel = 78;
			9407: Pixel = 79;
			9408: Pixel = 90;
			9409: Pixel = 82;
			9410: Pixel = 57;
			9411: Pixel = 66;
			9412: Pixel = 57;
			9413: Pixel = 57;
			9414: Pixel = 59;
			9415: Pixel = 56;
			9416: Pixel = 54;
			9417: Pixel = 60;
			9418: Pixel = 60;
			9419: Pixel = 58;
			9420: Pixel = 55;
			9421: Pixel = 56;
			9422: Pixel = 56;
			9423: Pixel = 52;
			9424: Pixel = 51;
			9425: Pixel = 50;
			9426: Pixel = 52;
			9427: Pixel = 36;
			9428: Pixel = 19;
			9429: Pixel = 22;
			9430: Pixel = 19;
			9431: Pixel = 40;
			9432: Pixel = 41;
			9433: Pixel = 28;
			9434: Pixel = 59;
			9435: Pixel = 48;
			9436: Pixel = 40;
			9437: Pixel = 36;
			9438: Pixel = 30;
			9439: Pixel = 39;
			9440: Pixel = 34;
			9441: Pixel = 45;
			9442: Pixel = 70;
			9443: Pixel = 93;
			9444: Pixel = 121;
			9445: Pixel = 99;
			9446: Pixel = 117;
			9447: Pixel = 134;
			9448: Pixel = 119;
			9449: Pixel = 93;
			9450: Pixel = 59;
			9451: Pixel = 45;
			9452: Pixel = 68;
			9453: Pixel = 82;
			9454: Pixel = 77;
			9455: Pixel = 76;
			9456: Pixel = 81;
			9457: Pixel = 84;
			9458: Pixel = 81;
			9459: Pixel = 83;
			9460: Pixel = 83;
			9461: Pixel = 80;
			9462: Pixel = 70;
			9463: Pixel = 81;
			9464: Pixel = 110;
			9465: Pixel = 117;
			9466: Pixel = 57;
			9467: Pixel = 34;
			9468: Pixel = 38;
			9469: Pixel = 40;
			9470: Pixel = 43;
			9471: Pixel = 47;
			9472: Pixel = 66;
			9473: Pixel = 51;
			9474: Pixel = 44;
			9475: Pixel = 51;
			9476: Pixel = 51;
			9477: Pixel = 59;
			9478: Pixel = 69;
			9479: Pixel = 81;
			9480: Pixel = 81;
			9481: Pixel = 71;
			9482: Pixel = 74;
			9483: Pixel = 68;
			9484: Pixel = 64;
			9485: Pixel = 57;
			9486: Pixel = 48;
			9487: Pixel = 50;
			9488: Pixel = 50;
			9489: Pixel = 66;
			9490: Pixel = 73;
			9491: Pixel = 90;
			9492: Pixel = 72;
			9493: Pixel = 138;
			9494: Pixel = 90;
			9495: Pixel = 137;
			9496: Pixel = 201;
			9497: Pixel = 243;
			9498: Pixel = 249;
			9499: Pixel = 247;
			9500: Pixel = 124;
			9501: Pixel = 104;
			9502: Pixel = 84;
			9503: Pixel = 75;
			9504: Pixel = 92;
			9505: Pixel = 81;
			9506: Pixel = 68;
			9507: Pixel = 78;
			9508: Pixel = 87;
			9509: Pixel = 75;
			9510: Pixel = 54;
			9511: Pixel = 64;
			9512: Pixel = 55;
			9513: Pixel = 55;
			9514: Pixel = 58;
			9515: Pixel = 55;
			9516: Pixel = 52;
			9517: Pixel = 58;
			9518: Pixel = 58;
			9519: Pixel = 57;
			9520: Pixel = 56;
			9521: Pixel = 57;
			9522: Pixel = 59;
			9523: Pixel = 53;
			9524: Pixel = 52;
			9525: Pixel = 48;
			9526: Pixel = 50;
			9527: Pixel = 39;
			9528: Pixel = 21;
			9529: Pixel = 18;
			9530: Pixel = 15;
			9531: Pixel = 38;
			9532: Pixel = 48;
			9533: Pixel = 45;
			9534: Pixel = 77;
			9535: Pixel = 35;
			9536: Pixel = 28;
			9537: Pixel = 36;
			9538: Pixel = 30;
			9539: Pixel = 50;
			9540: Pixel = 44;
			9541: Pixel = 45;
			9542: Pixel = 63;
			9543: Pixel = 96;
			9544: Pixel = 153;
			9545: Pixel = 97;
			9546: Pixel = 113;
			9547: Pixel = 136;
			9548: Pixel = 131;
			9549: Pixel = 104;
			9550: Pixel = 74;
			9551: Pixel = 42;
			9552: Pixel = 56;
			9553: Pixel = 78;
			9554: Pixel = 81;
			9555: Pixel = 75;
			9556: Pixel = 81;
			9557: Pixel = 83;
			9558: Pixel = 79;
			9559: Pixel = 81;
			9560: Pixel = 80;
			9561: Pixel = 76;
			9562: Pixel = 80;
			9563: Pixel = 95;
			9564: Pixel = 108;
			9565: Pixel = 117;
			9566: Pixel = 54;
			9567: Pixel = 33;
			9568: Pixel = 36;
			9569: Pixel = 38;
			9570: Pixel = 42;
			9571: Pixel = 51;
			9572: Pixel = 65;
			9573: Pixel = 53;
			9574: Pixel = 50;
			9575: Pixel = 54;
			9576: Pixel = 57;
			9577: Pixel = 67;
			9578: Pixel = 73;
			9579: Pixel = 71;
			9580: Pixel = 69;
			9581: Pixel = 76;
			9582: Pixel = 84;
			9583: Pixel = 91;
			9584: Pixel = 82;
			9585: Pixel = 74;
			9586: Pixel = 54;
			9587: Pixel = 53;
			9588: Pixel = 53;
			9589: Pixel = 70;
			9590: Pixel = 67;
			9591: Pixel = 89;
			9592: Pixel = 79;
			9593: Pixel = 115;
			9594: Pixel = 170;
			9595: Pixel = 221;
			9596: Pixel = 246;
			9597: Pixel = 248;
			9598: Pixel = 245;
			9599: Pixel = 220;
			9600: Pixel = 114;
			9601: Pixel = 111;
			9602: Pixel = 95;
			9603: Pixel = 70;
			9604: Pixel = 84;
			9605: Pixel = 78;
			9606: Pixel = 68;
			9607: Pixel = 75;
			9608: Pixel = 86;
			9609: Pixel = 76;
			9610: Pixel = 52;
			9611: Pixel = 60;
			9612: Pixel = 56;
			9613: Pixel = 51;
			9614: Pixel = 56;
			9615: Pixel = 55;
			9616: Pixel = 53;
			9617: Pixel = 54;
			9618: Pixel = 55;
			9619: Pixel = 55;
			9620: Pixel = 54;
			9621: Pixel = 53;
			9622: Pixel = 59;
			9623: Pixel = 51;
			9624: Pixel = 50;
			9625: Pixel = 49;
			9626: Pixel = 49;
			9627: Pixel = 47;
			9628: Pixel = 21;
			9629: Pixel = 50;
			9630: Pixel = 72;
			9631: Pixel = 73;
			9632: Pixel = 69;
			9633: Pixel = 45;
			9634: Pixel = 51;
			9635: Pixel = 24;
			9636: Pixel = 23;
			9637: Pixel = 31;
			9638: Pixel = 33;
			9639: Pixel = 46;
			9640: Pixel = 43;
			9641: Pixel = 37;
			9642: Pixel = 56;
			9643: Pixel = 98;
			9644: Pixel = 177;
			9645: Pixel = 95;
			9646: Pixel = 111;
			9647: Pixel = 138;
			9648: Pixel = 146;
			9649: Pixel = 116;
			9650: Pixel = 87;
			9651: Pixel = 45;
			9652: Pixel = 48;
			9653: Pixel = 68;
			9654: Pixel = 69;
			9655: Pixel = 67;
			9656: Pixel = 72;
			9657: Pixel = 74;
			9658: Pixel = 71;
			9659: Pixel = 70;
			9660: Pixel = 85;
			9661: Pixel = 99;
			9662: Pixel = 111;
			9663: Pixel = 109;
			9664: Pixel = 105;
			9665: Pixel = 116;
			9666: Pixel = 55;
			9667: Pixel = 37;
			9668: Pixel = 37;
			9669: Pixel = 38;
			9670: Pixel = 41;
			9671: Pixel = 54;
			9672: Pixel = 64;
			9673: Pixel = 47;
			9674: Pixel = 58;
			9675: Pixel = 67;
			9676: Pixel = 67;
			9677: Pixel = 81;
			9678: Pixel = 62;
			9679: Pixel = 67;
			9680: Pixel = 73;
			9681: Pixel = 87;
			9682: Pixel = 104;
			9683: Pixel = 108;
			9684: Pixel = 88;
			9685: Pixel = 82;
			9686: Pixel = 67;
			9687: Pixel = 55;
			9688: Pixel = 58;
			9689: Pixel = 77;
			9690: Pixel = 71;
			9691: Pixel = 81;
			9692: Pixel = 126;
			9693: Pixel = 180;
			9694: Pixel = 235;
			9695: Pixel = 248;
			9696: Pixel = 248;
			9697: Pixel = 245;
			9698: Pixel = 209;
			9699: Pixel = 150;
			9700: Pixel = 100;
			9701: Pixel = 117;
			9702: Pixel = 103;
			9703: Pixel = 68;
			9704: Pixel = 76;
			9705: Pixel = 76;
			9706: Pixel = 70;
			9707: Pixel = 72;
			9708: Pixel = 83;
			9709: Pixel = 68;
			9710: Pixel = 54;
			9711: Pixel = 56;
			9712: Pixel = 56;
			9713: Pixel = 48;
			9714: Pixel = 49;
			9715: Pixel = 53;
			9716: Pixel = 49;
			9717: Pixel = 50;
			9718: Pixel = 53;
			9719: Pixel = 53;
			9720: Pixel = 51;
			9721: Pixel = 49;
			9722: Pixel = 58;
			9723: Pixel = 54;
			9724: Pixel = 49;
			9725: Pixel = 46;
			9726: Pixel = 51;
			9727: Pixel = 41;
			9728: Pixel = 44;
			9729: Pixel = 122;
			9730: Pixel = 104;
			9731: Pixel = 92;
			9732: Pixel = 76;
			9733: Pixel = 43;
			9734: Pixel = 39;
			9735: Pixel = 26;
			9736: Pixel = 22;
			9737: Pixel = 30;
			9738: Pixel = 36;
			9739: Pixel = 40;
			9740: Pixel = 38;
			9741: Pixel = 32;
			9742: Pixel = 50;
			9743: Pixel = 95;
			9744: Pixel = 185;
			9745: Pixel = 98;
			9746: Pixel = 114;
			9747: Pixel = 136;
			9748: Pixel = 162;
			9749: Pixel = 128;
			9750: Pixel = 97;
			9751: Pixel = 62;
			9752: Pixel = 53;
			9753: Pixel = 53;
			9754: Pixel = 62;
			9755: Pixel = 61;
			9756: Pixel = 61;
			9757: Pixel = 74;
			9758: Pixel = 80;
			9759: Pixel = 79;
			9760: Pixel = 100;
			9761: Pixel = 122;
			9762: Pixel = 134;
			9763: Pixel = 114;
			9764: Pixel = 101;
			9765: Pixel = 122;
			9766: Pixel = 71;
			9767: Pixel = 37;
			9768: Pixel = 40;
			9769: Pixel = 41;
			9770: Pixel = 57;
			9771: Pixel = 71;
			9772: Pixel = 59;
			9773: Pixel = 72;
			9774: Pixel = 82;
			9775: Pixel = 87;
			9776: Pixel = 98;
			9777: Pixel = 106;
			9778: Pixel = 64;
			9779: Pixel = 70;
			9780: Pixel = 94;
			9781: Pixel = 107;
			9782: Pixel = 118;
			9783: Pixel = 105;
			9784: Pixel = 92;
			9785: Pixel = 89;
			9786: Pixel = 83;
			9787: Pixel = 65;
			9788: Pixel = 58;
			9789: Pixel = 85;
			9790: Pixel = 96;
			9791: Pixel = 145;
			9792: Pixel = 203;
			9793: Pixel = 242;
			9794: Pixel = 247;
			9795: Pixel = 249;
			9796: Pixel = 241;
			9797: Pixel = 196;
			9798: Pixel = 131;
			9799: Pixel = 84;
			9800: Pixel = 115;
			9801: Pixel = 123;
			9802: Pixel = 116;
			9803: Pixel = 81;
			9804: Pixel = 77;
			9805: Pixel = 78;
			9806: Pixel = 73;
			9807: Pixel = 72;
			9808: Pixel = 78;
			9809: Pixel = 64;
			9810: Pixel = 51;
			9811: Pixel = 54;
			9812: Pixel = 57;
			9813: Pixel = 50;
			9814: Pixel = 47;
			9815: Pixel = 54;
			9816: Pixel = 49;
			9817: Pixel = 46;
			9818: Pixel = 55;
			9819: Pixel = 54;
			9820: Pixel = 51;
			9821: Pixel = 50;
			9822: Pixel = 53;
			9823: Pixel = 46;
			9824: Pixel = 43;
			9825: Pixel = 30;
			9826: Pixel = 35;
			9827: Pixel = 36;
			9828: Pixel = 52;
			9829: Pixel = 93;
			9830: Pixel = 76;
			9831: Pixel = 73;
			9832: Pixel = 77;
			9833: Pixel = 54;
			9834: Pixel = 39;
			9835: Pixel = 27;
			9836: Pixel = 23;
			9837: Pixel = 29;
			9838: Pixel = 36;
			9839: Pixel = 35;
			9840: Pixel = 38;
			9841: Pixel = 40;
			9842: Pixel = 45;
			9843: Pixel = 87;
			9844: Pixel = 180;
			9845: Pixel = 102;
			9846: Pixel = 112;
			9847: Pixel = 133;
			9848: Pixel = 164;
			9849: Pixel = 141;
			9850: Pixel = 107;
			9851: Pixel = 76;
			9852: Pixel = 60;
			9853: Pixel = 61;
			9854: Pixel = 56;
			9855: Pixel = 75;
			9856: Pixel = 98;
			9857: Pixel = 95;
			9858: Pixel = 109;
			9859: Pixel = 121;
			9860: Pixel = 121;
			9861: Pixel = 122;
			9862: Pixel = 131;
			9863: Pixel = 116;
			9864: Pixel = 101;
			9865: Pixel = 128;
			9866: Pixel = 120;
			9867: Pixel = 38;
			9868: Pixel = 44;
			9869: Pixel = 43;
			9870: Pixel = 56;
			9871: Pixel = 70;
			9872: Pixel = 54;
			9873: Pixel = 73;
			9874: Pixel = 63;
			9875: Pixel = 111;
			9876: Pixel = 152;
			9877: Pixel = 175;
			9878: Pixel = 79;
			9879: Pixel = 85;
			9880: Pixel = 105;
			9881: Pixel = 106;
			9882: Pixel = 120;
			9883: Pixel = 113;
			9884: Pixel = 106;
			9885: Pixel = 92;
			9886: Pixel = 90;
			9887: Pixel = 85;
			9888: Pixel = 73;
			9889: Pixel = 119;
			9890: Pixel = 178;
			9891: Pixel = 224;
			9892: Pixel = 245;
			9893: Pixel = 247;
			9894: Pixel = 248;
			9895: Pixel = 229;
			9896: Pixel = 182;
			9897: Pixel = 116;
			9898: Pixel = 80;
			9899: Pixel = 78;
			9900: Pixel = 156;
			9901: Pixel = 139;
			9902: Pixel = 133;
			9903: Pixel = 95;
			9904: Pixel = 76;
			9905: Pixel = 77;
			9906: Pixel = 72;
			9907: Pixel = 73;
			9908: Pixel = 83;
			9909: Pixel = 66;
			9910: Pixel = 50;
			9911: Pixel = 54;
			9912: Pixel = 58;
			9913: Pixel = 54;
			9914: Pixel = 44;
			9915: Pixel = 52;
			9916: Pixel = 50;
			9917: Pixel = 43;
			9918: Pixel = 55;
			9919: Pixel = 54;
			9920: Pixel = 49;
			9921: Pixel = 55;
			9922: Pixel = 42;
			9923: Pixel = 32;
			9924: Pixel = 35;
			9925: Pixel = 27;
			9926: Pixel = 29;
			9927: Pixel = 39;
			9928: Pixel = 39;
			9929: Pixel = 81;
			9930: Pixel = 86;
			9931: Pixel = 74;
			9932: Pixel = 68;
			9933: Pixel = 68;
			9934: Pixel = 39;
			9935: Pixel = 28;
			9936: Pixel = 23;
			9937: Pixel = 27;
			9938: Pixel = 40;
			9939: Pixel = 45;
			9940: Pixel = 47;
			9941: Pixel = 46;
			9942: Pixel = 46;
			9943: Pixel = 77;
			9944: Pixel = 150;
			9945: Pixel = 103;
			9946: Pixel = 111;
			9947: Pixel = 133;
			9948: Pixel = 166;
			9949: Pixel = 155;
			9950: Pixel = 118;
			9951: Pixel = 86;
			9952: Pixel = 60;
			9953: Pixel = 60;
			9954: Pixel = 84;
			9955: Pixel = 127;
			9956: Pixel = 105;
			9957: Pixel = 88;
			9958: Pixel = 118;
			9959: Pixel = 128;
			9960: Pixel = 133;
			9961: Pixel = 137;
			9962: Pixel = 131;
			9963: Pixel = 109;
			9964: Pixel = 105;
			9965: Pixel = 124;
			9966: Pixel = 156;
			9967: Pixel = 57;
			9968: Pixel = 41;
			9969: Pixel = 44;
			9970: Pixel = 43;
			9971: Pixel = 51;
			9972: Pixel = 47;
			9973: Pixel = 47;
			9974: Pixel = 50;
			9975: Pixel = 112;
			9976: Pixel = 180;
			9977: Pixel = 156;
			9978: Pixel = 91;
			9979: Pixel = 96;
			9980: Pixel = 93;
			9981: Pixel = 106;
			9982: Pixel = 118;
			9983: Pixel = 118;
			9984: Pixel = 115;
			9985: Pixel = 93;
			9986: Pixel = 88;
			9987: Pixel = 104;
			9988: Pixel = 136;
			9989: Pixel = 198;
			9990: Pixel = 236;
			9991: Pixel = 248;
			9992: Pixel = 246;
			9993: Pixel = 243;
			9994: Pixel = 214;
			9995: Pixel = 174;
			9996: Pixel = 124;
			9997: Pixel = 78;
			9998: Pixel = 79;
			9999: Pixel = 80;
		endcase
	end
endmodule