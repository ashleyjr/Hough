module InHandle(
	input wire			nReset,                                                      // Common to all
	input wire			Clk,                                                        // Common to all
	output reg	[7:0]	Pixel,
	output reg			Frame,
	output reg			Line
);

	parameter COLS = 150;
	parameter ROWS = 150;
	
	reg [7:0] col;
	reg [7:0] row;
	
	always @ (posedge Clk or negedge nReset) begin
		if(!nReset) begin   
			Frame <= 0;
	    	Line  <= 0;							
			row <= ROWS-1;
			col <= COLS-1;						// Zero on first pixel	
		end else begin
			if(col == (COLS-1)) begin			// Get ready for next column
	    		Line <= 1;
				col <= 0;
				row <= row + 1;
				if(row == (ROWS-1)) begin		// Get ready for next row
					Frame <= 1;
					row <= 0;
				end
			end else begin
				Line <= 0;
				Frame <= 0;
				col = col + 1;
			end
		end
	end

	always @ (*) begin
		case(col + (row*COLS))


			0: Pixel = 162;
			1: Pixel = 160;
			2: Pixel = 161;
			3: Pixel = 159;
			4: Pixel = 157;
			5: Pixel = 158;
			6: Pixel = 155;
			7: Pixel = 155;
			8: Pixel = 154;
			9: Pixel = 155;
			10: Pixel = 159;
			11: Pixel = 164;
			12: Pixel = 168;
			13: Pixel = 173;
			14: Pixel = 171;
			15: Pixel = 167;
			16: Pixel = 155;
			17: Pixel = 139;
			18: Pixel = 108;
			19: Pixel = 92;
			20: Pixel = 96;
			21: Pixel = 102;
			22: Pixel = 104;
			23: Pixel = 108;
			24: Pixel = 106;
			25: Pixel = 108;
			26: Pixel = 108;
			27: Pixel = 108;
			28: Pixel = 109;
			29: Pixel = 105;
			30: Pixel = 108;
			31: Pixel = 114;
			32: Pixel = 117;
			33: Pixel = 120;
			34: Pixel = 122;
			35: Pixel = 126;
			36: Pixel = 126;
			37: Pixel = 131;
			38: Pixel = 130;
			39: Pixel = 130;
			40: Pixel = 134;
			41: Pixel = 130;
			42: Pixel = 129;
			43: Pixel = 129;
			44: Pixel = 129;
			45: Pixel = 130;
			46: Pixel = 133;
			47: Pixel = 131;
			48: Pixel = 133;
			49: Pixel = 133;
			50: Pixel = 133;
			51: Pixel = 134;
			52: Pixel = 133;
			53: Pixel = 131;
			54: Pixel = 134;
			55: Pixel = 132;
			56: Pixel = 133;
			57: Pixel = 134;
			58: Pixel = 135;
			59: Pixel = 134;
			60: Pixel = 134;
			61: Pixel = 135;
			62: Pixel = 132;
			63: Pixel = 130;
			64: Pixel = 131;
			65: Pixel = 130;
			66: Pixel = 132;
			67: Pixel = 132;
			68: Pixel = 131;
			69: Pixel = 130;
			70: Pixel = 133;
			71: Pixel = 133;
			72: Pixel = 135;
			73: Pixel = 131;
			74: Pixel = 133;
			75: Pixel = 138;
			76: Pixel = 129;
			77: Pixel = 130;
			78: Pixel = 132;
			79: Pixel = 129;
			80: Pixel = 128;
			81: Pixel = 132;
			82: Pixel = 129;
			83: Pixel = 129;
			84: Pixel = 129;
			85: Pixel = 130;
			86: Pixel = 128;
			87: Pixel = 126;
			88: Pixel = 127;
			89: Pixel = 123;
			90: Pixel = 121;
			91: Pixel = 117;
			92: Pixel = 111;
			93: Pixel = 103;
			94: Pixel = 114;
			95: Pixel = 132;
			96: Pixel = 143;
			97: Pixel = 151;
			98: Pixel = 157;
			99: Pixel = 161;
			100: Pixel = 154;
			101: Pixel = 150;
			102: Pixel = 151;
			103: Pixel = 154;
			104: Pixel = 154;
			105: Pixel = 156;
			106: Pixel = 155;
			107: Pixel = 153;
			108: Pixel = 153;
			109: Pixel = 152;
			110: Pixel = 152;
			111: Pixel = 154;
			112: Pixel = 153;
			113: Pixel = 157;
			114: Pixel = 155;
			115: Pixel = 158;
			116: Pixel = 156;
			117: Pixel = 153;
			118: Pixel = 188;
			119: Pixel = 210;
			120: Pixel = 214;
			121: Pixel = 218;
			122: Pixel = 214;
			123: Pixel = 168;
			124: Pixel = 105;
			125: Pixel = 103;
			126: Pixel = 113;
			127: Pixel = 118;
			128: Pixel = 121;
			129: Pixel = 121;
			130: Pixel = 120;
			131: Pixel = 122;
			132: Pixel = 123;
			133: Pixel = 120;
			134: Pixel = 122;
			135: Pixel = 121;
			136: Pixel = 123;
			137: Pixel = 124;
			138: Pixel = 125;
			139: Pixel = 123;
			140: Pixel = 121;
			141: Pixel = 126;
			142: Pixel = 125;
			143: Pixel = 124;
			144: Pixel = 124;
			145: Pixel = 118;
			146: Pixel = 115;
			147: Pixel = 127;
			148: Pixel = 174;
			149: Pixel = 161;
			150: Pixel = 161;
			151: Pixel = 159;
			152: Pixel = 160;
			153: Pixel = 157;
			154: Pixel = 155;
			155: Pixel = 156;
			156: Pixel = 153;
			157: Pixel = 155;
			158: Pixel = 153;
			159: Pixel = 155;
			160: Pixel = 157;
			161: Pixel = 164;
			162: Pixel = 169;
			163: Pixel = 172;
			164: Pixel = 171;
			165: Pixel = 167;
			166: Pixel = 153;
			167: Pixel = 134;
			168: Pixel = 108;
			169: Pixel = 92;
			170: Pixel = 95;
			171: Pixel = 100;
			172: Pixel = 105;
			173: Pixel = 107;
			174: Pixel = 105;
			175: Pixel = 106;
			176: Pixel = 106;
			177: Pixel = 106;
			178: Pixel = 107;
			179: Pixel = 105;
			180: Pixel = 108;
			181: Pixel = 113;
			182: Pixel = 118;
			183: Pixel = 121;
			184: Pixel = 123;
			185: Pixel = 125;
			186: Pixel = 125;
			187: Pixel = 129;
			188: Pixel = 131;
			189: Pixel = 130;
			190: Pixel = 132;
			191: Pixel = 130;
			192: Pixel = 129;
			193: Pixel = 130;
			194: Pixel = 129;
			195: Pixel = 131;
			196: Pixel = 132;
			197: Pixel = 132;
			198: Pixel = 134;
			199: Pixel = 133;
			200: Pixel = 133;
			201: Pixel = 134;
			202: Pixel = 132;
			203: Pixel = 131;
			204: Pixel = 132;
			205: Pixel = 131;
			206: Pixel = 133;
			207: Pixel = 133;
			208: Pixel = 134;
			209: Pixel = 133;
			210: Pixel = 133;
			211: Pixel = 135;
			212: Pixel = 132;
			213: Pixel = 129;
			214: Pixel = 131;
			215: Pixel = 130;
			216: Pixel = 132;
			217: Pixel = 132;
			218: Pixel = 129;
			219: Pixel = 130;
			220: Pixel = 133;
			221: Pixel = 133;
			222: Pixel = 133;
			223: Pixel = 131;
			224: Pixel = 132;
			225: Pixel = 136;
			226: Pixel = 130;
			227: Pixel = 129;
			228: Pixel = 130;
			229: Pixel = 129;
			230: Pixel = 128;
			231: Pixel = 130;
			232: Pixel = 127;
			233: Pixel = 129;
			234: Pixel = 129;
			235: Pixel = 129;
			236: Pixel = 128;
			237: Pixel = 127;
			238: Pixel = 126;
			239: Pixel = 122;
			240: Pixel = 121;
			241: Pixel = 117;
			242: Pixel = 111;
			243: Pixel = 102;
			244: Pixel = 113;
			245: Pixel = 130;
			246: Pixel = 142;
			247: Pixel = 151;
			248: Pixel = 157;
			249: Pixel = 160;
			250: Pixel = 155;
			251: Pixel = 151;
			252: Pixel = 151;
			253: Pixel = 152;
			254: Pixel = 153;
			255: Pixel = 154;
			256: Pixel = 155;
			257: Pixel = 153;
			258: Pixel = 152;
			259: Pixel = 152;
			260: Pixel = 153;
			261: Pixel = 154;
			262: Pixel = 153;
			263: Pixel = 155;
			264: Pixel = 155;
			265: Pixel = 157;
			266: Pixel = 156;
			267: Pixel = 151;
			268: Pixel = 183;
			269: Pixel = 209;
			270: Pixel = 214;
			271: Pixel = 218;
			272: Pixel = 216;
			273: Pixel = 178;
			274: Pixel = 109;
			275: Pixel = 101;
			276: Pixel = 113;
			277: Pixel = 118;
			278: Pixel = 120;
			279: Pixel = 121;
			280: Pixel = 120;
			281: Pixel = 123;
			282: Pixel = 123;
			283: Pixel = 120;
			284: Pixel = 121;
			285: Pixel = 122;
			286: Pixel = 124;
			287: Pixel = 124;
			288: Pixel = 124;
			289: Pixel = 123;
			290: Pixel = 121;
			291: Pixel = 125;
			292: Pixel = 125;
			293: Pixel = 125;
			294: Pixel = 125;
			295: Pixel = 118;
			296: Pixel = 118;
			297: Pixel = 131;
			298: Pixel = 151;
			299: Pixel = 120;
			300: Pixel = 156;
			301: Pixel = 157;
			302: Pixel = 157;
			303: Pixel = 156;
			304: Pixel = 154;
			305: Pixel = 155;
			306: Pixel = 154;
			307: Pixel = 153;
			308: Pixel = 153;
			309: Pixel = 153;
			310: Pixel = 156;
			311: Pixel = 165;
			312: Pixel = 170;
			313: Pixel = 171;
			314: Pixel = 171;
			315: Pixel = 164;
			316: Pixel = 149;
			317: Pixel = 130;
			318: Pixel = 108;
			319: Pixel = 89;
			320: Pixel = 90;
			321: Pixel = 97;
			322: Pixel = 102;
			323: Pixel = 104;
			324: Pixel = 102;
			325: Pixel = 104;
			326: Pixel = 104;
			327: Pixel = 104;
			328: Pixel = 104;
			329: Pixel = 105;
			330: Pixel = 108;
			331: Pixel = 111;
			332: Pixel = 116;
			333: Pixel = 121;
			334: Pixel = 124;
			335: Pixel = 124;
			336: Pixel = 124;
			337: Pixel = 127;
			338: Pixel = 128;
			339: Pixel = 129;
			340: Pixel = 129;
			341: Pixel = 129;
			342: Pixel = 130;
			343: Pixel = 131;
			344: Pixel = 129;
			345: Pixel = 130;
			346: Pixel = 130;
			347: Pixel = 131;
			348: Pixel = 133;
			349: Pixel = 133;
			350: Pixel = 133;
			351: Pixel = 132;
			352: Pixel = 133;
			353: Pixel = 131;
			354: Pixel = 132;
			355: Pixel = 132;
			356: Pixel = 133;
			357: Pixel = 131;
			358: Pixel = 131;
			359: Pixel = 130;
			360: Pixel = 129;
			361: Pixel = 131;
			362: Pixel = 132;
			363: Pixel = 130;
			364: Pixel = 127;
			365: Pixel = 128;
			366: Pixel = 132;
			367: Pixel = 131;
			368: Pixel = 127;
			369: Pixel = 129;
			370: Pixel = 130;
			371: Pixel = 131;
			372: Pixel = 130;
			373: Pixel = 130;
			374: Pixel = 130;
			375: Pixel = 132;
			376: Pixel = 131;
			377: Pixel = 128;
			378: Pixel = 128;
			379: Pixel = 128;
			380: Pixel = 127;
			381: Pixel = 127;
			382: Pixel = 126;
			383: Pixel = 127;
			384: Pixel = 128;
			385: Pixel = 128;
			386: Pixel = 127;
			387: Pixel = 126;
			388: Pixel = 125;
			389: Pixel = 123;
			390: Pixel = 120;
			391: Pixel = 116;
			392: Pixel = 111;
			393: Pixel = 105;
			394: Pixel = 106;
			395: Pixel = 121;
			396: Pixel = 136;
			397: Pixel = 147;
			398: Pixel = 153;
			399: Pixel = 159;
			400: Pixel = 158;
			401: Pixel = 153;
			402: Pixel = 152;
			403: Pixel = 153;
			404: Pixel = 154;
			405: Pixel = 153;
			406: Pixel = 154;
			407: Pixel = 155;
			408: Pixel = 154;
			409: Pixel = 153;
			410: Pixel = 154;
			411: Pixel = 153;
			412: Pixel = 153;
			413: Pixel = 154;
			414: Pixel = 154;
			415: Pixel = 154;
			416: Pixel = 153;
			417: Pixel = 150;
			418: Pixel = 159;
			419: Pixel = 198;
			420: Pixel = 212;
			421: Pixel = 215;
			422: Pixel = 218;
			423: Pixel = 207;
			424: Pixel = 144;
			425: Pixel = 100;
			426: Pixel = 109;
			427: Pixel = 114;
			428: Pixel = 118;
			429: Pixel = 119;
			430: Pixel = 120;
			431: Pixel = 121;
			432: Pixel = 122;
			433: Pixel = 120;
			434: Pixel = 120;
			435: Pixel = 123;
			436: Pixel = 124;
			437: Pixel = 123;
			438: Pixel = 122;
			439: Pixel = 124;
			440: Pixel = 123;
			441: Pixel = 124;
			442: Pixel = 126;
			443: Pixel = 125;
			444: Pixel = 127;
			445: Pixel = 126;
			446: Pixel = 128;
			447: Pixel = 108;
			448: Pixel = 61;
			449: Pixel = 44;
			450: Pixel = 157;
			451: Pixel = 155;
			452: Pixel = 155;
			453: Pixel = 156;
			454: Pixel = 156;
			455: Pixel = 156;
			456: Pixel = 155;
			457: Pixel = 153;
			458: Pixel = 154;
			459: Pixel = 154;
			460: Pixel = 161;
			461: Pixel = 167;
			462: Pixel = 169;
			463: Pixel = 169;
			464: Pixel = 168;
			465: Pixel = 163;
			466: Pixel = 146;
			467: Pixel = 130;
			468: Pixel = 106;
			469: Pixel = 89;
			470: Pixel = 91;
			471: Pixel = 96;
			472: Pixel = 100;
			473: Pixel = 103;
			474: Pixel = 105;
			475: Pixel = 107;
			476: Pixel = 105;
			477: Pixel = 102;
			478: Pixel = 103;
			479: Pixel = 102;
			480: Pixel = 109;
			481: Pixel = 112;
			482: Pixel = 116;
			483: Pixel = 120;
			484: Pixel = 122;
			485: Pixel = 123;
			486: Pixel = 125;
			487: Pixel = 126;
			488: Pixel = 127;
			489: Pixel = 128;
			490: Pixel = 128;
			491: Pixel = 130;
			492: Pixel = 132;
			493: Pixel = 130;
			494: Pixel = 129;
			495: Pixel = 129;
			496: Pixel = 130;
			497: Pixel = 130;
			498: Pixel = 132;
			499: Pixel = 131;
			500: Pixel = 133;
			501: Pixel = 133;
			502: Pixel = 131;
			503: Pixel = 131;
			504: Pixel = 132;
			505: Pixel = 132;
			506: Pixel = 131;
			507: Pixel = 130;
			508: Pixel = 131;
			509: Pixel = 131;
			510: Pixel = 130;
			511: Pixel = 131;
			512: Pixel = 130;
			513: Pixel = 129;
			514: Pixel = 129;
			515: Pixel = 129;
			516: Pixel = 129;
			517: Pixel = 130;
			518: Pixel = 128;
			519: Pixel = 129;
			520: Pixel = 131;
			521: Pixel = 133;
			522: Pixel = 131;
			523: Pixel = 130;
			524: Pixel = 129;
			525: Pixel = 129;
			526: Pixel = 130;
			527: Pixel = 131;
			528: Pixel = 130;
			529: Pixel = 128;
			530: Pixel = 129;
			531: Pixel = 128;
			532: Pixel = 127;
			533: Pixel = 128;
			534: Pixel = 126;
			535: Pixel = 127;
			536: Pixel = 128;
			537: Pixel = 127;
			538: Pixel = 127;
			539: Pixel = 123;
			540: Pixel = 120;
			541: Pixel = 117;
			542: Pixel = 112;
			543: Pixel = 109;
			544: Pixel = 104;
			545: Pixel = 109;
			546: Pixel = 130;
			547: Pixel = 142;
			548: Pixel = 151;
			549: Pixel = 157;
			550: Pixel = 159;
			551: Pixel = 156;
			552: Pixel = 155;
			553: Pixel = 156;
			554: Pixel = 158;
			555: Pixel = 159;
			556: Pixel = 158;
			557: Pixel = 157;
			558: Pixel = 156;
			559: Pixel = 153;
			560: Pixel = 155;
			561: Pixel = 155;
			562: Pixel = 153;
			563: Pixel = 152;
			564: Pixel = 151;
			565: Pixel = 153;
			566: Pixel = 153;
			567: Pixel = 153;
			568: Pixel = 148;
			569: Pixel = 175;
			570: Pixel = 207;
			571: Pixel = 214;
			572: Pixel = 217;
			573: Pixel = 218;
			574: Pixel = 188;
			575: Pixel = 117;
			576: Pixel = 102;
			577: Pixel = 111;
			578: Pixel = 115;
			579: Pixel = 119;
			580: Pixel = 119;
			581: Pixel = 121;
			582: Pixel = 121;
			583: Pixel = 120;
			584: Pixel = 118;
			585: Pixel = 121;
			586: Pixel = 121;
			587: Pixel = 121;
			588: Pixel = 123;
			589: Pixel = 123;
			590: Pixel = 123;
			591: Pixel = 125;
			592: Pixel = 125;
			593: Pixel = 124;
			594: Pixel = 131;
			595: Pixel = 134;
			596: Pixel = 104;
			597: Pixel = 59;
			598: Pixel = 42;
			599: Pixel = 48;
			600: Pixel = 157;
			601: Pixel = 156;
			602: Pixel = 155;
			603: Pixel = 156;
			604: Pixel = 155;
			605: Pixel = 155;
			606: Pixel = 155;
			607: Pixel = 153;
			608: Pixel = 155;
			609: Pixel = 160;
			610: Pixel = 166;
			611: Pixel = 167;
			612: Pixel = 168;
			613: Pixel = 167;
			614: Pixel = 165;
			615: Pixel = 159;
			616: Pixel = 146;
			617: Pixel = 128;
			618: Pixel = 106;
			619: Pixel = 90;
			620: Pixel = 90;
			621: Pixel = 97;
			622: Pixel = 102;
			623: Pixel = 104;
			624: Pixel = 107;
			625: Pixel = 106;
			626: Pixel = 104;
			627: Pixel = 104;
			628: Pixel = 103;
			629: Pixel = 101;
			630: Pixel = 108;
			631: Pixel = 112;
			632: Pixel = 116;
			633: Pixel = 119;
			634: Pixel = 123;
			635: Pixel = 124;
			636: Pixel = 125;
			637: Pixel = 127;
			638: Pixel = 127;
			639: Pixel = 128;
			640: Pixel = 128;
			641: Pixel = 131;
			642: Pixel = 131;
			643: Pixel = 130;
			644: Pixel = 130;
			645: Pixel = 129;
			646: Pixel = 130;
			647: Pixel = 132;
			648: Pixel = 132;
			649: Pixel = 131;
			650: Pixel = 134;
			651: Pixel = 133;
			652: Pixel = 131;
			653: Pixel = 132;
			654: Pixel = 133;
			655: Pixel = 132;
			656: Pixel = 129;
			657: Pixel = 132;
			658: Pixel = 132;
			659: Pixel = 131;
			660: Pixel = 132;
			661: Pixel = 132;
			662: Pixel = 132;
			663: Pixel = 131;
			664: Pixel = 130;
			665: Pixel = 129;
			666: Pixel = 131;
			667: Pixel = 130;
			668: Pixel = 129;
			669: Pixel = 130;
			670: Pixel = 133;
			671: Pixel = 135;
			672: Pixel = 133;
			673: Pixel = 131;
			674: Pixel = 131;
			675: Pixel = 130;
			676: Pixel = 130;
			677: Pixel = 129;
			678: Pixel = 130;
			679: Pixel = 128;
			680: Pixel = 129;
			681: Pixel = 126;
			682: Pixel = 127;
			683: Pixel = 128;
			684: Pixel = 128;
			685: Pixel = 128;
			686: Pixel = 128;
			687: Pixel = 128;
			688: Pixel = 128;
			689: Pixel = 125;
			690: Pixel = 122;
			691: Pixel = 117;
			692: Pixel = 113;
			693: Pixel = 114;
			694: Pixel = 107;
			695: Pixel = 104;
			696: Pixel = 120;
			697: Pixel = 140;
			698: Pixel = 148;
			699: Pixel = 154;
			700: Pixel = 159;
			701: Pixel = 161;
			702: Pixel = 160;
			703: Pixel = 158;
			704: Pixel = 161;
			705: Pixel = 161;
			706: Pixel = 162;
			707: Pixel = 158;
			708: Pixel = 157;
			709: Pixel = 157;
			710: Pixel = 155;
			711: Pixel = 153;
			712: Pixel = 154;
			713: Pixel = 154;
			714: Pixel = 151;
			715: Pixel = 151;
			716: Pixel = 152;
			717: Pixel = 152;
			718: Pixel = 149;
			719: Pixel = 153;
			720: Pixel = 193;
			721: Pixel = 212;
			722: Pixel = 217;
			723: Pixel = 219;
			724: Pixel = 213;
			725: Pixel = 161;
			726: Pixel = 105;
			727: Pixel = 107;
			728: Pixel = 112;
			729: Pixel = 117;
			730: Pixel = 117;
			731: Pixel = 119;
			732: Pixel = 121;
			733: Pixel = 121;
			734: Pixel = 120;
			735: Pixel = 122;
			736: Pixel = 121;
			737: Pixel = 123;
			738: Pixel = 123;
			739: Pixel = 125;
			740: Pixel = 125;
			741: Pixel = 126;
			742: Pixel = 127;
			743: Pixel = 132;
			744: Pixel = 133;
			745: Pixel = 97;
			746: Pixel = 53;
			747: Pixel = 47;
			748: Pixel = 48;
			749: Pixel = 49;
			750: Pixel = 156;
			751: Pixel = 156;
			752: Pixel = 155;
			753: Pixel = 157;
			754: Pixel = 157;
			755: Pixel = 157;
			756: Pixel = 155;
			757: Pixel = 153;
			758: Pixel = 157;
			759: Pixel = 163;
			760: Pixel = 165;
			761: Pixel = 166;
			762: Pixel = 166;
			763: Pixel = 164;
			764: Pixel = 163;
			765: Pixel = 157;
			766: Pixel = 146;
			767: Pixel = 132;
			768: Pixel = 109;
			769: Pixel = 90;
			770: Pixel = 90;
			771: Pixel = 97;
			772: Pixel = 101;
			773: Pixel = 103;
			774: Pixel = 106;
			775: Pixel = 106;
			776: Pixel = 104;
			777: Pixel = 104;
			778: Pixel = 103;
			779: Pixel = 102;
			780: Pixel = 107;
			781: Pixel = 113;
			782: Pixel = 116;
			783: Pixel = 119;
			784: Pixel = 121;
			785: Pixel = 124;
			786: Pixel = 123;
			787: Pixel = 127;
			788: Pixel = 128;
			789: Pixel = 129;
			790: Pixel = 129;
			791: Pixel = 131;
			792: Pixel = 130;
			793: Pixel = 131;
			794: Pixel = 132;
			795: Pixel = 130;
			796: Pixel = 130;
			797: Pixel = 131;
			798: Pixel = 132;
			799: Pixel = 130;
			800: Pixel = 132;
			801: Pixel = 133;
			802: Pixel = 133;
			803: Pixel = 131;
			804: Pixel = 131;
			805: Pixel = 132;
			806: Pixel = 130;
			807: Pixel = 131;
			808: Pixel = 134;
			809: Pixel = 131;
			810: Pixel = 133;
			811: Pixel = 131;
			812: Pixel = 131;
			813: Pixel = 133;
			814: Pixel = 131;
			815: Pixel = 129;
			816: Pixel = 131;
			817: Pixel = 131;
			818: Pixel = 128;
			819: Pixel = 129;
			820: Pixel = 132;
			821: Pixel = 134;
			822: Pixel = 136;
			823: Pixel = 132;
			824: Pixel = 131;
			825: Pixel = 131;
			826: Pixel = 130;
			827: Pixel = 133;
			828: Pixel = 128;
			829: Pixel = 127;
			830: Pixel = 129;
			831: Pixel = 130;
			832: Pixel = 127;
			833: Pixel = 126;
			834: Pixel = 128;
			835: Pixel = 130;
			836: Pixel = 129;
			837: Pixel = 126;
			838: Pixel = 128;
			839: Pixel = 126;
			840: Pixel = 123;
			841: Pixel = 120;
			842: Pixel = 115;
			843: Pixel = 113;
			844: Pixel = 108;
			845: Pixel = 103;
			846: Pixel = 112;
			847: Pixel = 133;
			848: Pixel = 145;
			849: Pixel = 153;
			850: Pixel = 158;
			851: Pixel = 162;
			852: Pixel = 162;
			853: Pixel = 160;
			854: Pixel = 160;
			855: Pixel = 163;
			856: Pixel = 162;
			857: Pixel = 161;
			858: Pixel = 158;
			859: Pixel = 159;
			860: Pixel = 158;
			861: Pixel = 155;
			862: Pixel = 153;
			863: Pixel = 155;
			864: Pixel = 152;
			865: Pixel = 151;
			866: Pixel = 152;
			867: Pixel = 151;
			868: Pixel = 151;
			869: Pixel = 146;
			870: Pixel = 167;
			871: Pixel = 205;
			872: Pixel = 215;
			873: Pixel = 218;
			874: Pixel = 219;
			875: Pixel = 199;
			876: Pixel = 129;
			877: Pixel = 100;
			878: Pixel = 110;
			879: Pixel = 114;
			880: Pixel = 116;
			881: Pixel = 119;
			882: Pixel = 123;
			883: Pixel = 122;
			884: Pixel = 123;
			885: Pixel = 122;
			886: Pixel = 123;
			887: Pixel = 124;
			888: Pixel = 125;
			889: Pixel = 127;
			890: Pixel = 128;
			891: Pixel = 131;
			892: Pixel = 134;
			893: Pixel = 133;
			894: Pixel = 94;
			895: Pixel = 47;
			896: Pixel = 46;
			897: Pixel = 48;
			898: Pixel = 48;
			899: Pixel = 46;
			900: Pixel = 156;
			901: Pixel = 155;
			902: Pixel = 156;
			903: Pixel = 157;
			904: Pixel = 158;
			905: Pixel = 157;
			906: Pixel = 155;
			907: Pixel = 154;
			908: Pixel = 158;
			909: Pixel = 165;
			910: Pixel = 166;
			911: Pixel = 164;
			912: Pixel = 164;
			913: Pixel = 162;
			914: Pixel = 160;
			915: Pixel = 158;
			916: Pixel = 147;
			917: Pixel = 134;
			918: Pixel = 111;
			919: Pixel = 90;
			920: Pixel = 92;
			921: Pixel = 97;
			922: Pixel = 101;
			923: Pixel = 108;
			924: Pixel = 104;
			925: Pixel = 103;
			926: Pixel = 104;
			927: Pixel = 102;
			928: Pixel = 103;
			929: Pixel = 103;
			930: Pixel = 107;
			931: Pixel = 112;
			932: Pixel = 114;
			933: Pixel = 119;
			934: Pixel = 120;
			935: Pixel = 123;
			936: Pixel = 124;
			937: Pixel = 125;
			938: Pixel = 127;
			939: Pixel = 129;
			940: Pixel = 130;
			941: Pixel = 129;
			942: Pixel = 129;
			943: Pixel = 130;
			944: Pixel = 129;
			945: Pixel = 129;
			946: Pixel = 130;
			947: Pixel = 130;
			948: Pixel = 131;
			949: Pixel = 130;
			950: Pixel = 132;
			951: Pixel = 132;
			952: Pixel = 129;
			953: Pixel = 130;
			954: Pixel = 129;
			955: Pixel = 130;
			956: Pixel = 130;
			957: Pixel = 131;
			958: Pixel = 131;
			959: Pixel = 128;
			960: Pixel = 131;
			961: Pixel = 130;
			962: Pixel = 128;
			963: Pixel = 129;
			964: Pixel = 129;
			965: Pixel = 130;
			966: Pixel = 130;
			967: Pixel = 129;
			968: Pixel = 127;
			969: Pixel = 128;
			970: Pixel = 131;
			971: Pixel = 132;
			972: Pixel = 135;
			973: Pixel = 132;
			974: Pixel = 130;
			975: Pixel = 130;
			976: Pixel = 130;
			977: Pixel = 131;
			978: Pixel = 129;
			979: Pixel = 128;
			980: Pixel = 128;
			981: Pixel = 126;
			982: Pixel = 126;
			983: Pixel = 125;
			984: Pixel = 127;
			985: Pixel = 127;
			986: Pixel = 127;
			987: Pixel = 126;
			988: Pixel = 128;
			989: Pixel = 124;
			990: Pixel = 123;
			991: Pixel = 123;
			992: Pixel = 117;
			993: Pixel = 111;
			994: Pixel = 109;
			995: Pixel = 105;
			996: Pixel = 108;
			997: Pixel = 126;
			998: Pixel = 144;
			999: Pixel = 152;
			1000: Pixel = 157;
			1001: Pixel = 162;
			1002: Pixel = 163;
			1003: Pixel = 161;
			1004: Pixel = 160;
			1005: Pixel = 160;
			1006: Pixel = 161;
			1007: Pixel = 160;
			1008: Pixel = 160;
			1009: Pixel = 155;
			1010: Pixel = 156;
			1011: Pixel = 155;
			1012: Pixel = 154;
			1013: Pixel = 152;
			1014: Pixel = 151;
			1015: Pixel = 151;
			1016: Pixel = 151;
			1017: Pixel = 150;
			1018: Pixel = 151;
			1019: Pixel = 148;
			1020: Pixel = 146;
			1021: Pixel = 186;
			1022: Pixel = 211;
			1023: Pixel = 216;
			1024: Pixel = 219;
			1025: Pixel = 217;
			1026: Pixel = 173;
			1027: Pixel = 107;
			1028: Pixel = 108;
			1029: Pixel = 112;
			1030: Pixel = 116;
			1031: Pixel = 118;
			1032: Pixel = 118;
			1033: Pixel = 122;
			1034: Pixel = 121;
			1035: Pixel = 121;
			1036: Pixel = 120;
			1037: Pixel = 126;
			1038: Pixel = 129;
			1039: Pixel = 129;
			1040: Pixel = 131;
			1041: Pixel = 135;
			1042: Pixel = 137;
			1043: Pixel = 94;
			1044: Pixel = 51;
			1045: Pixel = 45;
			1046: Pixel = 52;
			1047: Pixel = 49;
			1048: Pixel = 47;
			1049: Pixel = 51;
			1050: Pixel = 154;
			1051: Pixel = 155;
			1052: Pixel = 158;
			1053: Pixel = 158;
			1054: Pixel = 157;
			1055: Pixel = 157;
			1056: Pixel = 156;
			1057: Pixel = 157;
			1058: Pixel = 163;
			1059: Pixel = 166;
			1060: Pixel = 167;
			1061: Pixel = 164;
			1062: Pixel = 162;
			1063: Pixel = 159;
			1064: Pixel = 160;
			1065: Pixel = 158;
			1066: Pixel = 148;
			1067: Pixel = 130;
			1068: Pixel = 105;
			1069: Pixel = 86;
			1070: Pixel = 88;
			1071: Pixel = 96;
			1072: Pixel = 101;
			1073: Pixel = 104;
			1074: Pixel = 104;
			1075: Pixel = 104;
			1076: Pixel = 105;
			1077: Pixel = 103;
			1078: Pixel = 102;
			1079: Pixel = 104;
			1080: Pixel = 108;
			1081: Pixel = 110;
			1082: Pixel = 114;
			1083: Pixel = 120;
			1084: Pixel = 120;
			1085: Pixel = 121;
			1086: Pixel = 124;
			1087: Pixel = 127;
			1088: Pixel = 128;
			1089: Pixel = 126;
			1090: Pixel = 129;
			1091: Pixel = 130;
			1092: Pixel = 128;
			1093: Pixel = 129;
			1094: Pixel = 129;
			1095: Pixel = 129;
			1096: Pixel = 129;
			1097: Pixel = 130;
			1098: Pixel = 129;
			1099: Pixel = 127;
			1100: Pixel = 131;
			1101: Pixel = 131;
			1102: Pixel = 130;
			1103: Pixel = 128;
			1104: Pixel = 130;
			1105: Pixel = 131;
			1106: Pixel = 134;
			1107: Pixel = 132;
			1108: Pixel = 129;
			1109: Pixel = 127;
			1110: Pixel = 126;
			1111: Pixel = 125;
			1112: Pixel = 125;
			1113: Pixel = 126;
			1114: Pixel = 126;
			1115: Pixel = 127;
			1116: Pixel = 126;
			1117: Pixel = 126;
			1118: Pixel = 127;
			1119: Pixel = 126;
			1120: Pixel = 128;
			1121: Pixel = 128;
			1122: Pixel = 130;
			1123: Pixel = 132;
			1124: Pixel = 130;
			1125: Pixel = 130;
			1126: Pixel = 132;
			1127: Pixel = 129;
			1128: Pixel = 127;
			1129: Pixel = 126;
			1130: Pixel = 128;
			1131: Pixel = 126;
			1132: Pixel = 126;
			1133: Pixel = 125;
			1134: Pixel = 127;
			1135: Pixel = 127;
			1136: Pixel = 125;
			1137: Pixel = 126;
			1138: Pixel = 127;
			1139: Pixel = 124;
			1140: Pixel = 123;
			1141: Pixel = 123;
			1142: Pixel = 118;
			1143: Pixel = 109;
			1144: Pixel = 108;
			1145: Pixel = 105;
			1146: Pixel = 112;
			1147: Pixel = 124;
			1148: Pixel = 140;
			1149: Pixel = 150;
			1150: Pixel = 158;
			1151: Pixel = 162;
			1152: Pixel = 161;
			1153: Pixel = 163;
			1154: Pixel = 160;
			1155: Pixel = 158;
			1156: Pixel = 159;
			1157: Pixel = 158;
			1158: Pixel = 159;
			1159: Pixel = 156;
			1160: Pixel = 155;
			1161: Pixel = 155;
			1162: Pixel = 155;
			1163: Pixel = 153;
			1164: Pixel = 152;
			1165: Pixel = 152;
			1166: Pixel = 151;
			1167: Pixel = 151;
			1168: Pixel = 150;
			1169: Pixel = 149;
			1170: Pixel = 143;
			1171: Pixel = 160;
			1172: Pixel = 202;
			1173: Pixel = 215;
			1174: Pixel = 218;
			1175: Pixel = 220;
			1176: Pixel = 208;
			1177: Pixel = 142;
			1178: Pixel = 100;
			1179: Pixel = 112;
			1180: Pixel = 115;
			1181: Pixel = 120;
			1182: Pixel = 121;
			1183: Pixel = 122;
			1184: Pixel = 122;
			1185: Pixel = 120;
			1186: Pixel = 120;
			1187: Pixel = 123;
			1188: Pixel = 124;
			1189: Pixel = 128;
			1190: Pixel = 135;
			1191: Pixel = 136;
			1192: Pixel = 91;
			1193: Pixel = 55;
			1194: Pixel = 49;
			1195: Pixel = 43;
			1196: Pixel = 44;
			1197: Pixel = 45;
			1198: Pixel = 51;
			1199: Pixel = 53;
			1200: Pixel = 157;
			1201: Pixel = 157;
			1202: Pixel = 157;
			1203: Pixel = 159;
			1204: Pixel = 158;
			1205: Pixel = 159;
			1206: Pixel = 158;
			1207: Pixel = 161;
			1208: Pixel = 167;
			1209: Pixel = 167;
			1210: Pixel = 166;
			1211: Pixel = 163;
			1212: Pixel = 158;
			1213: Pixel = 157;
			1214: Pixel = 161;
			1215: Pixel = 161;
			1216: Pixel = 149;
			1217: Pixel = 129;
			1218: Pixel = 104;
			1219: Pixel = 87;
			1220: Pixel = 86;
			1221: Pixel = 97;
			1222: Pixel = 101;
			1223: Pixel = 104;
			1224: Pixel = 105;
			1225: Pixel = 105;
			1226: Pixel = 104;
			1227: Pixel = 103;
			1228: Pixel = 103;
			1229: Pixel = 104;
			1230: Pixel = 107;
			1231: Pixel = 109;
			1232: Pixel = 115;
			1233: Pixel = 120;
			1234: Pixel = 121;
			1235: Pixel = 123;
			1236: Pixel = 124;
			1237: Pixel = 126;
			1238: Pixel = 126;
			1239: Pixel = 126;
			1240: Pixel = 127;
			1241: Pixel = 127;
			1242: Pixel = 127;
			1243: Pixel = 128;
			1244: Pixel = 129;
			1245: Pixel = 130;
			1246: Pixel = 129;
			1247: Pixel = 130;
			1248: Pixel = 130;
			1249: Pixel = 129;
			1250: Pixel = 128;
			1251: Pixel = 130;
			1252: Pixel = 129;
			1253: Pixel = 127;
			1254: Pixel = 129;
			1255: Pixel = 131;
			1256: Pixel = 134;
			1257: Pixel = 134;
			1258: Pixel = 130;
			1259: Pixel = 125;
			1260: Pixel = 124;
			1261: Pixel = 122;
			1262: Pixel = 123;
			1263: Pixel = 123;
			1264: Pixel = 128;
			1265: Pixel = 127;
			1266: Pixel = 124;
			1267: Pixel = 125;
			1268: Pixel = 125;
			1269: Pixel = 126;
			1270: Pixel = 127;
			1271: Pixel = 129;
			1272: Pixel = 128;
			1273: Pixel = 130;
			1274: Pixel = 130;
			1275: Pixel = 131;
			1276: Pixel = 132;
			1277: Pixel = 128;
			1278: Pixel = 126;
			1279: Pixel = 126;
			1280: Pixel = 127;
			1281: Pixel = 128;
			1282: Pixel = 127;
			1283: Pixel = 126;
			1284: Pixel = 126;
			1285: Pixel = 126;
			1286: Pixel = 125;
			1287: Pixel = 127;
			1288: Pixel = 128;
			1289: Pixel = 125;
			1290: Pixel = 122;
			1291: Pixel = 120;
			1292: Pixel = 119;
			1293: Pixel = 114;
			1294: Pixel = 110;
			1295: Pixel = 106;
			1296: Pixel = 113;
			1297: Pixel = 126;
			1298: Pixel = 138;
			1299: Pixel = 149;
			1300: Pixel = 157;
			1301: Pixel = 159;
			1302: Pixel = 161;
			1303: Pixel = 161;
			1304: Pixel = 159;
			1305: Pixel = 158;
			1306: Pixel = 159;
			1307: Pixel = 158;
			1308: Pixel = 158;
			1309: Pixel = 157;
			1310: Pixel = 156;
			1311: Pixel = 155;
			1312: Pixel = 157;
			1313: Pixel = 154;
			1314: Pixel = 154;
			1315: Pixel = 156;
			1316: Pixel = 153;
			1317: Pixel = 152;
			1318: Pixel = 151;
			1319: Pixel = 148;
			1320: Pixel = 146;
			1321: Pixel = 144;
			1322: Pixel = 182;
			1323: Pixel = 212;
			1324: Pixel = 216;
			1325: Pixel = 220;
			1326: Pixel = 220;
			1327: Pixel = 188;
			1328: Pixel = 112;
			1329: Pixel = 106;
			1330: Pixel = 114;
			1331: Pixel = 117;
			1332: Pixel = 121;
			1333: Pixel = 122;
			1334: Pixel = 121;
			1335: Pixel = 121;
			1336: Pixel = 121;
			1337: Pixel = 124;
			1338: Pixel = 126;
			1339: Pixel = 132;
			1340: Pixel = 134;
			1341: Pixel = 90;
			1342: Pixel = 44;
			1343: Pixel = 43;
			1344: Pixel = 46;
			1345: Pixel = 43;
			1346: Pixel = 47;
			1347: Pixel = 49;
			1348: Pixel = 50;
			1349: Pixel = 54;
			1350: Pixel = 158;
			1351: Pixel = 157;
			1352: Pixel = 157;
			1353: Pixel = 159;
			1354: Pixel = 160;
			1355: Pixel = 160;
			1356: Pixel = 162;
			1357: Pixel = 167;
			1358: Pixel = 168;
			1359: Pixel = 168;
			1360: Pixel = 167;
			1361: Pixel = 161;
			1362: Pixel = 158;
			1363: Pixel = 157;
			1364: Pixel = 161;
			1365: Pixel = 161;
			1366: Pixel = 150;
			1367: Pixel = 131;
			1368: Pixel = 105;
			1369: Pixel = 89;
			1370: Pixel = 91;
			1371: Pixel = 97;
			1372: Pixel = 99;
			1373: Pixel = 105;
			1374: Pixel = 107;
			1375: Pixel = 106;
			1376: Pixel = 104;
			1377: Pixel = 101;
			1378: Pixel = 102;
			1379: Pixel = 103;
			1380: Pixel = 106;
			1381: Pixel = 110;
			1382: Pixel = 114;
			1383: Pixel = 119;
			1384: Pixel = 122;
			1385: Pixel = 123;
			1386: Pixel = 122;
			1387: Pixel = 125;
			1388: Pixel = 127;
			1389: Pixel = 127;
			1390: Pixel = 128;
			1391: Pixel = 127;
			1392: Pixel = 126;
			1393: Pixel = 127;
			1394: Pixel = 128;
			1395: Pixel = 129;
			1396: Pixel = 129;
			1397: Pixel = 130;
			1398: Pixel = 130;
			1399: Pixel = 131;
			1400: Pixel = 131;
			1401: Pixel = 128;
			1402: Pixel = 130;
			1403: Pixel = 130;
			1404: Pixel = 128;
			1405: Pixel = 130;
			1406: Pixel = 131;
			1407: Pixel = 131;
			1408: Pixel = 129;
			1409: Pixel = 127;
			1410: Pixel = 124;
			1411: Pixel = 122;
			1412: Pixel = 121;
			1413: Pixel = 122;
			1414: Pixel = 122;
			1415: Pixel = 126;
			1416: Pixel = 125;
			1417: Pixel = 125;
			1418: Pixel = 124;
			1419: Pixel = 124;
			1420: Pixel = 125;
			1421: Pixel = 129;
			1422: Pixel = 129;
			1423: Pixel = 128;
			1424: Pixel = 129;
			1425: Pixel = 132;
			1426: Pixel = 130;
			1427: Pixel = 127;
			1428: Pixel = 127;
			1429: Pixel = 126;
			1430: Pixel = 128;
			1431: Pixel = 127;
			1432: Pixel = 127;
			1433: Pixel = 125;
			1434: Pixel = 127;
			1435: Pixel = 125;
			1436: Pixel = 126;
			1437: Pixel = 127;
			1438: Pixel = 127;
			1439: Pixel = 127;
			1440: Pixel = 124;
			1441: Pixel = 119;
			1442: Pixel = 117;
			1443: Pixel = 112;
			1444: Pixel = 110;
			1445: Pixel = 107;
			1446: Pixel = 112;
			1447: Pixel = 126;
			1448: Pixel = 136;
			1449: Pixel = 145;
			1450: Pixel = 153;
			1451: Pixel = 156;
			1452: Pixel = 159;
			1453: Pixel = 160;
			1454: Pixel = 158;
			1455: Pixel = 157;
			1456: Pixel = 159;
			1457: Pixel = 159;
			1458: Pixel = 158;
			1459: Pixel = 156;
			1460: Pixel = 156;
			1461: Pixel = 155;
			1462: Pixel = 156;
			1463: Pixel = 155;
			1464: Pixel = 156;
			1465: Pixel = 156;
			1466: Pixel = 154;
			1467: Pixel = 154;
			1468: Pixel = 152;
			1469: Pixel = 151;
			1470: Pixel = 148;
			1471: Pixel = 140;
			1472: Pixel = 151;
			1473: Pixel = 196;
			1474: Pixel = 211;
			1475: Pixel = 218;
			1476: Pixel = 221;
			1477: Pixel = 218;
			1478: Pixel = 164;
			1479: Pixel = 106;
			1480: Pixel = 110;
			1481: Pixel = 115;
			1482: Pixel = 117;
			1483: Pixel = 120;
			1484: Pixel = 121;
			1485: Pixel = 121;
			1486: Pixel = 124;
			1487: Pixel = 124;
			1488: Pixel = 131;
			1489: Pixel = 133;
			1490: Pixel = 95;
			1491: Pixel = 45;
			1492: Pixel = 42;
			1493: Pixel = 50;
			1494: Pixel = 47;
			1495: Pixel = 49;
			1496: Pixel = 51;
			1497: Pixel = 50;
			1498: Pixel = 49;
			1499: Pixel = 55;
			1500: Pixel = 158;
			1501: Pixel = 157;
			1502: Pixel = 159;
			1503: Pixel = 161;
			1504: Pixel = 161;
			1505: Pixel = 163;
			1506: Pixel = 166;
			1507: Pixel = 168;
			1508: Pixel = 168;
			1509: Pixel = 166;
			1510: Pixel = 165;
			1511: Pixel = 159;
			1512: Pixel = 158;
			1513: Pixel = 158;
			1514: Pixel = 160;
			1515: Pixel = 160;
			1516: Pixel = 146;
			1517: Pixel = 130;
			1518: Pixel = 104;
			1519: Pixel = 87;
			1520: Pixel = 89;
			1521: Pixel = 97;
			1522: Pixel = 100;
			1523: Pixel = 104;
			1524: Pixel = 103;
			1525: Pixel = 103;
			1526: Pixel = 103;
			1527: Pixel = 102;
			1528: Pixel = 101;
			1529: Pixel = 103;
			1530: Pixel = 106;
			1531: Pixel = 111;
			1532: Pixel = 115;
			1533: Pixel = 117;
			1534: Pixel = 120;
			1535: Pixel = 120;
			1536: Pixel = 123;
			1537: Pixel = 123;
			1538: Pixel = 126;
			1539: Pixel = 127;
			1540: Pixel = 126;
			1541: Pixel = 129;
			1542: Pixel = 127;
			1543: Pixel = 126;
			1544: Pixel = 125;
			1545: Pixel = 127;
			1546: Pixel = 130;
			1547: Pixel = 128;
			1548: Pixel = 128;
			1549: Pixel = 127;
			1550: Pixel = 128;
			1551: Pixel = 128;
			1552: Pixel = 130;
			1553: Pixel = 130;
			1554: Pixel = 129;
			1555: Pixel = 128;
			1556: Pixel = 130;
			1557: Pixel = 130;
			1558: Pixel = 125;
			1559: Pixel = 125;
			1560: Pixel = 124;
			1561: Pixel = 124;
			1562: Pixel = 121;
			1563: Pixel = 122;
			1564: Pixel = 124;
			1565: Pixel = 126;
			1566: Pixel = 126;
			1567: Pixel = 121;
			1568: Pixel = 121;
			1569: Pixel = 122;
			1570: Pixel = 123;
			1571: Pixel = 127;
			1572: Pixel = 128;
			1573: Pixel = 130;
			1574: Pixel = 129;
			1575: Pixel = 131;
			1576: Pixel = 131;
			1577: Pixel = 128;
			1578: Pixel = 127;
			1579: Pixel = 128;
			1580: Pixel = 128;
			1581: Pixel = 126;
			1582: Pixel = 126;
			1583: Pixel = 125;
			1584: Pixel = 125;
			1585: Pixel = 126;
			1586: Pixel = 125;
			1587: Pixel = 126;
			1588: Pixel = 126;
			1589: Pixel = 126;
			1590: Pixel = 123;
			1591: Pixel = 120;
			1592: Pixel = 117;
			1593: Pixel = 114;
			1594: Pixel = 112;
			1595: Pixel = 107;
			1596: Pixel = 112;
			1597: Pixel = 122;
			1598: Pixel = 135;
			1599: Pixel = 142;
			1600: Pixel = 150;
			1601: Pixel = 154;
			1602: Pixel = 156;
			1603: Pixel = 158;
			1604: Pixel = 158;
			1605: Pixel = 156;
			1606: Pixel = 157;
			1607: Pixel = 158;
			1608: Pixel = 157;
			1609: Pixel = 155;
			1610: Pixel = 158;
			1611: Pixel = 155;
			1612: Pixel = 157;
			1613: Pixel = 156;
			1614: Pixel = 155;
			1615: Pixel = 155;
			1616: Pixel = 155;
			1617: Pixel = 155;
			1618: Pixel = 151;
			1619: Pixel = 151;
			1620: Pixel = 149;
			1621: Pixel = 145;
			1622: Pixel = 140;
			1623: Pixel = 173;
			1624: Pixel = 210;
			1625: Pixel = 218;
			1626: Pixel = 221;
			1627: Pixel = 222;
			1628: Pixel = 203;
			1629: Pixel = 128;
			1630: Pixel = 99;
			1631: Pixel = 111;
			1632: Pixel = 115;
			1633: Pixel = 118;
			1634: Pixel = 123;
			1635: Pixel = 123;
			1636: Pixel = 126;
			1637: Pixel = 131;
			1638: Pixel = 132;
			1639: Pixel = 91;
			1640: Pixel = 44;
			1641: Pixel = 41;
			1642: Pixel = 45;
			1643: Pixel = 51;
			1644: Pixel = 54;
			1645: Pixel = 52;
			1646: Pixel = 52;
			1647: Pixel = 50;
			1648: Pixel = 52;
			1649: Pixel = 50;
			1650: Pixel = 161;
			1651: Pixel = 159;
			1652: Pixel = 160;
			1653: Pixel = 161;
			1654: Pixel = 162;
			1655: Pixel = 166;
			1656: Pixel = 168;
			1657: Pixel = 166;
			1658: Pixel = 164;
			1659: Pixel = 164;
			1660: Pixel = 162;
			1661: Pixel = 159;
			1662: Pixel = 158;
			1663: Pixel = 160;
			1664: Pixel = 161;
			1665: Pixel = 159;
			1666: Pixel = 147;
			1667: Pixel = 129;
			1668: Pixel = 102;
			1669: Pixel = 83;
			1670: Pixel = 86;
			1671: Pixel = 95;
			1672: Pixel = 101;
			1673: Pixel = 103;
			1674: Pixel = 102;
			1675: Pixel = 101;
			1676: Pixel = 102;
			1677: Pixel = 102;
			1678: Pixel = 103;
			1679: Pixel = 102;
			1680: Pixel = 105;
			1681: Pixel = 112;
			1682: Pixel = 115;
			1683: Pixel = 118;
			1684: Pixel = 120;
			1685: Pixel = 119;
			1686: Pixel = 121;
			1687: Pixel = 123;
			1688: Pixel = 124;
			1689: Pixel = 125;
			1690: Pixel = 124;
			1691: Pixel = 127;
			1692: Pixel = 125;
			1693: Pixel = 123;
			1694: Pixel = 124;
			1695: Pixel = 126;
			1696: Pixel = 128;
			1697: Pixel = 128;
			1698: Pixel = 128;
			1699: Pixel = 125;
			1700: Pixel = 127;
			1701: Pixel = 128;
			1702: Pixel = 130;
			1703: Pixel = 130;
			1704: Pixel = 128;
			1705: Pixel = 127;
			1706: Pixel = 129;
			1707: Pixel = 127;
			1708: Pixel = 127;
			1709: Pixel = 126;
			1710: Pixel = 126;
			1711: Pixel = 124;
			1712: Pixel = 122;
			1713: Pixel = 124;
			1714: Pixel = 121;
			1715: Pixel = 122;
			1716: Pixel = 120;
			1717: Pixel = 120;
			1718: Pixel = 120;
			1719: Pixel = 121;
			1720: Pixel = 123;
			1721: Pixel = 125;
			1722: Pixel = 127;
			1723: Pixel = 128;
			1724: Pixel = 130;
			1725: Pixel = 130;
			1726: Pixel = 129;
			1727: Pixel = 127;
			1728: Pixel = 126;
			1729: Pixel = 126;
			1730: Pixel = 128;
			1731: Pixel = 127;
			1732: Pixel = 126;
			1733: Pixel = 126;
			1734: Pixel = 125;
			1735: Pixel = 125;
			1736: Pixel = 126;
			1737: Pixel = 125;
			1738: Pixel = 126;
			1739: Pixel = 125;
			1740: Pixel = 123;
			1741: Pixel = 118;
			1742: Pixel = 117;
			1743: Pixel = 118;
			1744: Pixel = 113;
			1745: Pixel = 108;
			1746: Pixel = 111;
			1747: Pixel = 123;
			1748: Pixel = 134;
			1749: Pixel = 142;
			1750: Pixel = 147;
			1751: Pixel = 151;
			1752: Pixel = 154;
			1753: Pixel = 156;
			1754: Pixel = 157;
			1755: Pixel = 157;
			1756: Pixel = 156;
			1757: Pixel = 156;
			1758: Pixel = 155;
			1759: Pixel = 155;
			1760: Pixel = 156;
			1761: Pixel = 153;
			1762: Pixel = 154;
			1763: Pixel = 157;
			1764: Pixel = 156;
			1765: Pixel = 155;
			1766: Pixel = 154;
			1767: Pixel = 153;
			1768: Pixel = 150;
			1769: Pixel = 149;
			1770: Pixel = 148;
			1771: Pixel = 145;
			1772: Pixel = 140;
			1773: Pixel = 146;
			1774: Pixel = 195;
			1775: Pixel = 216;
			1776: Pixel = 220;
			1777: Pixel = 223;
			1778: Pixel = 221;
			1779: Pixel = 177;
			1780: Pixel = 103;
			1781: Pixel = 105;
			1782: Pixel = 111;
			1783: Pixel = 115;
			1784: Pixel = 118;
			1785: Pixel = 122;
			1786: Pixel = 129;
			1787: Pixel = 132;
			1788: Pixel = 90;
			1789: Pixel = 44;
			1790: Pixel = 43;
			1791: Pixel = 44;
			1792: Pixel = 47;
			1793: Pixel = 56;
			1794: Pixel = 57;
			1795: Pixel = 55;
			1796: Pixel = 51;
			1797: Pixel = 50;
			1798: Pixel = 47;
			1799: Pixel = 47;
			1800: Pixel = 160;
			1801: Pixel = 161;
			1802: Pixel = 159;
			1803: Pixel = 161;
			1804: Pixel = 165;
			1805: Pixel = 169;
			1806: Pixel = 165;
			1807: Pixel = 160;
			1808: Pixel = 159;
			1809: Pixel = 159;
			1810: Pixel = 158;
			1811: Pixel = 161;
			1812: Pixel = 158;
			1813: Pixel = 159;
			1814: Pixel = 160;
			1815: Pixel = 159;
			1816: Pixel = 147;
			1817: Pixel = 128;
			1818: Pixel = 101;
			1819: Pixel = 83;
			1820: Pixel = 87;
			1821: Pixel = 95;
			1822: Pixel = 102;
			1823: Pixel = 103;
			1824: Pixel = 102;
			1825: Pixel = 103;
			1826: Pixel = 103;
			1827: Pixel = 102;
			1828: Pixel = 101;
			1829: Pixel = 102;
			1830: Pixel = 105;
			1831: Pixel = 110;
			1832: Pixel = 115;
			1833: Pixel = 120;
			1834: Pixel = 119;
			1835: Pixel = 120;
			1836: Pixel = 123;
			1837: Pixel = 123;
			1838: Pixel = 123;
			1839: Pixel = 123;
			1840: Pixel = 126;
			1841: Pixel = 125;
			1842: Pixel = 124;
			1843: Pixel = 125;
			1844: Pixel = 127;
			1845: Pixel = 128;
			1846: Pixel = 128;
			1847: Pixel = 127;
			1848: Pixel = 126;
			1849: Pixel = 127;
			1850: Pixel = 128;
			1851: Pixel = 128;
			1852: Pixel = 128;
			1853: Pixel = 129;
			1854: Pixel = 128;
			1855: Pixel = 127;
			1856: Pixel = 129;
			1857: Pixel = 127;
			1858: Pixel = 127;
			1859: Pixel = 127;
			1860: Pixel = 128;
			1861: Pixel = 124;
			1862: Pixel = 123;
			1863: Pixel = 121;
			1864: Pixel = 119;
			1865: Pixel = 119;
			1866: Pixel = 120;
			1867: Pixel = 118;
			1868: Pixel = 115;
			1869: Pixel = 113;
			1870: Pixel = 115;
			1871: Pixel = 121;
			1872: Pixel = 125;
			1873: Pixel = 127;
			1874: Pixel = 129;
			1875: Pixel = 128;
			1876: Pixel = 126;
			1877: Pixel = 126;
			1878: Pixel = 127;
			1879: Pixel = 125;
			1880: Pixel = 127;
			1881: Pixel = 130;
			1882: Pixel = 126;
			1883: Pixel = 128;
			1884: Pixel = 127;
			1885: Pixel = 126;
			1886: Pixel = 125;
			1887: Pixel = 126;
			1888: Pixel = 127;
			1889: Pixel = 123;
			1890: Pixel = 122;
			1891: Pixel = 119;
			1892: Pixel = 115;
			1893: Pixel = 114;
			1894: Pixel = 114;
			1895: Pixel = 109;
			1896: Pixel = 112;
			1897: Pixel = 121;
			1898: Pixel = 132;
			1899: Pixel = 140;
			1900: Pixel = 145;
			1901: Pixel = 148;
			1902: Pixel = 152;
			1903: Pixel = 153;
			1904: Pixel = 155;
			1905: Pixel = 157;
			1906: Pixel = 155;
			1907: Pixel = 154;
			1908: Pixel = 154;
			1909: Pixel = 154;
			1910: Pixel = 153;
			1911: Pixel = 153;
			1912: Pixel = 153;
			1913: Pixel = 154;
			1914: Pixel = 156;
			1915: Pixel = 154;
			1916: Pixel = 152;
			1917: Pixel = 149;
			1918: Pixel = 147;
			1919: Pixel = 146;
			1920: Pixel = 145;
			1921: Pixel = 143;
			1922: Pixel = 141;
			1923: Pixel = 138;
			1924: Pixel = 169;
			1925: Pixel = 210;
			1926: Pixel = 218;
			1927: Pixel = 221;
			1928: Pixel = 223;
			1929: Pixel = 210;
			1930: Pixel = 138;
			1931: Pixel = 98;
			1932: Pixel = 108;
			1933: Pixel = 111;
			1934: Pixel = 113;
			1935: Pixel = 123;
			1936: Pixel = 131;
			1937: Pixel = 93;
			1938: Pixel = 47;
			1939: Pixel = 42;
			1940: Pixel = 45;
			1941: Pixel = 47;
			1942: Pixel = 52;
			1943: Pixel = 58;
			1944: Pixel = 55;
			1945: Pixel = 52;
			1946: Pixel = 51;
			1947: Pixel = 46;
			1948: Pixel = 45;
			1949: Pixel = 44;
			1950: Pixel = 161;
			1951: Pixel = 161;
			1952: Pixel = 159;
			1953: Pixel = 162;
			1954: Pixel = 168;
			1955: Pixel = 166;
			1956: Pixel = 157;
			1957: Pixel = 154;
			1958: Pixel = 153;
			1959: Pixel = 153;
			1960: Pixel = 157;
			1961: Pixel = 163;
			1962: Pixel = 160;
			1963: Pixel = 159;
			1964: Pixel = 162;
			1965: Pixel = 159;
			1966: Pixel = 149;
			1967: Pixel = 131;
			1968: Pixel = 103;
			1969: Pixel = 84;
			1970: Pixel = 87;
			1971: Pixel = 95;
			1972: Pixel = 99;
			1973: Pixel = 103;
			1974: Pixel = 105;
			1975: Pixel = 104;
			1976: Pixel = 103;
			1977: Pixel = 103;
			1978: Pixel = 102;
			1979: Pixel = 103;
			1980: Pixel = 108;
			1981: Pixel = 111;
			1982: Pixel = 115;
			1983: Pixel = 119;
			1984: Pixel = 120;
			1985: Pixel = 122;
			1986: Pixel = 123;
			1987: Pixel = 123;
			1988: Pixel = 124;
			1989: Pixel = 125;
			1990: Pixel = 126;
			1991: Pixel = 125;
			1992: Pixel = 125;
			1993: Pixel = 127;
			1994: Pixel = 128;
			1995: Pixel = 128;
			1996: Pixel = 129;
			1997: Pixel = 128;
			1998: Pixel = 124;
			1999: Pixel = 129;
			2000: Pixel = 131;
			2001: Pixel = 128;
			2002: Pixel = 131;
			2003: Pixel = 128;
			2004: Pixel = 127;
			2005: Pixel = 126;
			2006: Pixel = 129;
			2007: Pixel = 129;
			2008: Pixel = 124;
			2009: Pixel = 124;
			2010: Pixel = 129;
			2011: Pixel = 134;
			2012: Pixel = 131;
			2013: Pixel = 133;
			2014: Pixel = 149;
			2015: Pixel = 161;
			2016: Pixel = 161;
			2017: Pixel = 158;
			2018: Pixel = 157;
			2019: Pixel = 151;
			2020: Pixel = 138;
			2021: Pixel = 123;
			2022: Pixel = 116;
			2023: Pixel = 114;
			2024: Pixel = 119;
			2025: Pixel = 123;
			2026: Pixel = 125;
			2027: Pixel = 126;
			2028: Pixel = 125;
			2029: Pixel = 127;
			2030: Pixel = 129;
			2031: Pixel = 129;
			2032: Pixel = 129;
			2033: Pixel = 127;
			2034: Pixel = 126;
			2035: Pixel = 127;
			2036: Pixel = 126;
			2037: Pixel = 126;
			2038: Pixel = 126;
			2039: Pixel = 125;
			2040: Pixel = 123;
			2041: Pixel = 119;
			2042: Pixel = 115;
			2043: Pixel = 115;
			2044: Pixel = 112;
			2045: Pixel = 107;
			2046: Pixel = 110;
			2047: Pixel = 119;
			2048: Pixel = 132;
			2049: Pixel = 139;
			2050: Pixel = 144;
			2051: Pixel = 145;
			2052: Pixel = 149;
			2053: Pixel = 150;
			2054: Pixel = 153;
			2055: Pixel = 155;
			2056: Pixel = 155;
			2057: Pixel = 153;
			2058: Pixel = 152;
			2059: Pixel = 153;
			2060: Pixel = 153;
			2061: Pixel = 154;
			2062: Pixel = 155;
			2063: Pixel = 153;
			2064: Pixel = 153;
			2065: Pixel = 152;
			2066: Pixel = 149;
			2067: Pixel = 148;
			2068: Pixel = 145;
			2069: Pixel = 144;
			2070: Pixel = 143;
			2071: Pixel = 143;
			2072: Pixel = 143;
			2073: Pixel = 141;
			2074: Pixel = 145;
			2075: Pixel = 191;
			2076: Pixel = 215;
			2077: Pixel = 220;
			2078: Pixel = 223;
			2079: Pixel = 221;
			2080: Pixel = 184;
			2081: Pixel = 109;
			2082: Pixel = 106;
			2083: Pixel = 112;
			2084: Pixel = 118;
			2085: Pixel = 125;
			2086: Pixel = 91;
			2087: Pixel = 47;
			2088: Pixel = 44;
			2089: Pixel = 46;
			2090: Pixel = 46;
			2091: Pixel = 50;
			2092: Pixel = 55;
			2093: Pixel = 59;
			2094: Pixel = 56;
			2095: Pixel = 52;
			2096: Pixel = 51;
			2097: Pixel = 45;
			2098: Pixel = 46;
			2099: Pixel = 47;
			2100: Pixel = 162;
			2101: Pixel = 160;
			2102: Pixel = 158;
			2103: Pixel = 166;
			2104: Pixel = 170;
			2105: Pixel = 162;
			2106: Pixel = 152;
			2107: Pixel = 147;
			2108: Pixel = 145;
			2109: Pixel = 147;
			2110: Pixel = 159;
			2111: Pixel = 163;
			2112: Pixel = 160;
			2113: Pixel = 160;
			2114: Pixel = 163;
			2115: Pixel = 159;
			2116: Pixel = 149;
			2117: Pixel = 132;
			2118: Pixel = 105;
			2119: Pixel = 86;
			2120: Pixel = 87;
			2121: Pixel = 94;
			2122: Pixel = 98;
			2123: Pixel = 103;
			2124: Pixel = 104;
			2125: Pixel = 105;
			2126: Pixel = 101;
			2127: Pixel = 104;
			2128: Pixel = 102;
			2129: Pixel = 103;
			2130: Pixel = 110;
			2131: Pixel = 112;
			2132: Pixel = 112;
			2133: Pixel = 119;
			2134: Pixel = 121;
			2135: Pixel = 121;
			2136: Pixel = 124;
			2137: Pixel = 125;
			2138: Pixel = 124;
			2139: Pixel = 126;
			2140: Pixel = 126;
			2141: Pixel = 126;
			2142: Pixel = 126;
			2143: Pixel = 129;
			2144: Pixel = 128;
			2145: Pixel = 128;
			2146: Pixel = 129;
			2147: Pixel = 127;
			2148: Pixel = 127;
			2149: Pixel = 127;
			2150: Pixel = 128;
			2151: Pixel = 132;
			2152: Pixel = 130;
			2153: Pixel = 128;
			2154: Pixel = 127;
			2155: Pixel = 124;
			2156: Pixel = 127;
			2157: Pixel = 138;
			2158: Pixel = 141;
			2159: Pixel = 144;
			2160: Pixel = 148;
			2161: Pixel = 146;
			2162: Pixel = 154;
			2163: Pixel = 165;
			2164: Pixel = 166;
			2165: Pixel = 176;
			2166: Pixel = 178;
			2167: Pixel = 178;
			2168: Pixel = 185;
			2169: Pixel = 186;
			2170: Pixel = 184;
			2171: Pixel = 179;
			2172: Pixel = 167;
			2173: Pixel = 142;
			2174: Pixel = 122;
			2175: Pixel = 113;
			2176: Pixel = 117;
			2177: Pixel = 123;
			2178: Pixel = 123;
			2179: Pixel = 125;
			2180: Pixel = 130;
			2181: Pixel = 130;
			2182: Pixel = 130;
			2183: Pixel = 127;
			2184: Pixel = 126;
			2185: Pixel = 125;
			2186: Pixel = 126;
			2187: Pixel = 126;
			2188: Pixel = 125;
			2189: Pixel = 125;
			2190: Pixel = 120;
			2191: Pixel = 119;
			2192: Pixel = 117;
			2193: Pixel = 112;
			2194: Pixel = 112;
			2195: Pixel = 108;
			2196: Pixel = 109;
			2197: Pixel = 119;
			2198: Pixel = 131;
			2199: Pixel = 140;
			2200: Pixel = 144;
			2201: Pixel = 143;
			2202: Pixel = 145;
			2203: Pixel = 148;
			2204: Pixel = 151;
			2205: Pixel = 154;
			2206: Pixel = 154;
			2207: Pixel = 154;
			2208: Pixel = 151;
			2209: Pixel = 153;
			2210: Pixel = 152;
			2211: Pixel = 153;
			2212: Pixel = 154;
			2213: Pixel = 153;
			2214: Pixel = 150;
			2215: Pixel = 150;
			2216: Pixel = 148;
			2217: Pixel = 145;
			2218: Pixel = 143;
			2219: Pixel = 144;
			2220: Pixel = 142;
			2221: Pixel = 142;
			2222: Pixel = 141;
			2223: Pixel = 141;
			2224: Pixel = 140;
			2225: Pixel = 163;
			2226: Pixel = 206;
			2227: Pixel = 217;
			2228: Pixel = 221;
			2229: Pixel = 224;
			2230: Pixel = 216;
			2231: Pixel = 153;
			2232: Pixel = 104;
			2233: Pixel = 116;
			2234: Pixel = 123;
			2235: Pixel = 90;
			2236: Pixel = 43;
			2237: Pixel = 41;
			2238: Pixel = 45;
			2239: Pixel = 44;
			2240: Pixel = 49;
			2241: Pixel = 54;
			2242: Pixel = 55;
			2243: Pixel = 58;
			2244: Pixel = 56;
			2245: Pixel = 50;
			2246: Pixel = 41;
			2247: Pixel = 45;
			2248: Pixel = 46;
			2249: Pixel = 47;
			2250: Pixel = 160;
			2251: Pixel = 159;
			2252: Pixel = 162;
			2253: Pixel = 168;
			2254: Pixel = 168;
			2255: Pixel = 158;
			2256: Pixel = 146;
			2257: Pixel = 138;
			2258: Pixel = 137;
			2259: Pixel = 144;
			2260: Pixel = 160;
			2261: Pixel = 164;
			2262: Pixel = 161;
			2263: Pixel = 161;
			2264: Pixel = 163;
			2265: Pixel = 160;
			2266: Pixel = 148;
			2267: Pixel = 131;
			2268: Pixel = 103;
			2269: Pixel = 83;
			2270: Pixel = 87;
			2271: Pixel = 93;
			2272: Pixel = 97;
			2273: Pixel = 103;
			2274: Pixel = 104;
			2275: Pixel = 102;
			2276: Pixel = 103;
			2277: Pixel = 103;
			2278: Pixel = 104;
			2279: Pixel = 105;
			2280: Pixel = 109;
			2281: Pixel = 113;
			2282: Pixel = 117;
			2283: Pixel = 120;
			2284: Pixel = 122;
			2285: Pixel = 120;
			2286: Pixel = 122;
			2287: Pixel = 126;
			2288: Pixel = 126;
			2289: Pixel = 124;
			2290: Pixel = 124;
			2291: Pixel = 126;
			2292: Pixel = 129;
			2293: Pixel = 129;
			2294: Pixel = 127;
			2295: Pixel = 129;
			2296: Pixel = 129;
			2297: Pixel = 129;
			2298: Pixel = 127;
			2299: Pixel = 127;
			2300: Pixel = 127;
			2301: Pixel = 127;
			2302: Pixel = 126;
			2303: Pixel = 127;
			2304: Pixel = 126;
			2305: Pixel = 134;
			2306: Pixel = 142;
			2307: Pixel = 149;
			2308: Pixel = 150;
			2309: Pixel = 142;
			2310: Pixel = 146;
			2311: Pixel = 150;
			2312: Pixel = 167;
			2313: Pixel = 167;
			2314: Pixel = 166;
			2315: Pixel = 176;
			2316: Pixel = 181;
			2317: Pixel = 178;
			2318: Pixel = 174;
			2319: Pixel = 168;
			2320: Pixel = 176;
			2321: Pixel = 184;
			2322: Pixel = 189;
			2323: Pixel = 193;
			2324: Pixel = 184;
			2325: Pixel = 161;
			2326: Pixel = 128;
			2327: Pixel = 110;
			2328: Pixel = 117;
			2329: Pixel = 123;
			2330: Pixel = 125;
			2331: Pixel = 126;
			2332: Pixel = 126;
			2333: Pixel = 127;
			2334: Pixel = 126;
			2335: Pixel = 124;
			2336: Pixel = 125;
			2337: Pixel = 124;
			2338: Pixel = 125;
			2339: Pixel = 121;
			2340: Pixel = 120;
			2341: Pixel = 118;
			2342: Pixel = 115;
			2343: Pixel = 113;
			2344: Pixel = 112;
			2345: Pixel = 106;
			2346: Pixel = 108;
			2347: Pixel = 118;
			2348: Pixel = 133;
			2349: Pixel = 140;
			2350: Pixel = 145;
			2351: Pixel = 143;
			2352: Pixel = 144;
			2353: Pixel = 146;
			2354: Pixel = 148;
			2355: Pixel = 152;
			2356: Pixel = 153;
			2357: Pixel = 153;
			2358: Pixel = 152;
			2359: Pixel = 151;
			2360: Pixel = 152;
			2361: Pixel = 150;
			2362: Pixel = 150;
			2363: Pixel = 150;
			2364: Pixel = 149;
			2365: Pixel = 146;
			2366: Pixel = 144;
			2367: Pixel = 144;
			2368: Pixel = 141;
			2369: Pixel = 141;
			2370: Pixel = 139;
			2371: Pixel = 140;
			2372: Pixel = 141;
			2373: Pixel = 141;
			2374: Pixel = 140;
			2375: Pixel = 141;
			2376: Pixel = 181;
			2377: Pixel = 213;
			2378: Pixel = 219;
			2379: Pixel = 224;
			2380: Pixel = 226;
			2381: Pixel = 202;
			2382: Pixel = 129;
			2383: Pixel = 119;
			2384: Pixel = 96;
			2385: Pixel = 46;
			2386: Pixel = 40;
			2387: Pixel = 45;
			2388: Pixel = 46;
			2389: Pixel = 46;
			2390: Pixel = 51;
			2391: Pixel = 54;
			2392: Pixel = 51;
			2393: Pixel = 51;
			2394: Pixel = 49;
			2395: Pixel = 47;
			2396: Pixel = 47;
			2397: Pixel = 48;
			2398: Pixel = 45;
			2399: Pixel = 44;
			2400: Pixel = 159;
			2401: Pixel = 161;
			2402: Pixel = 168;
			2403: Pixel = 170;
			2404: Pixel = 162;
			2405: Pixel = 151;
			2406: Pixel = 137;
			2407: Pixel = 126;
			2408: Pixel = 131;
			2409: Pixel = 147;
			2410: Pixel = 160;
			2411: Pixel = 164;
			2412: Pixel = 163;
			2413: Pixel = 164;
			2414: Pixel = 165;
			2415: Pixel = 161;
			2416: Pixel = 149;
			2417: Pixel = 131;
			2418: Pixel = 101;
			2419: Pixel = 79;
			2420: Pixel = 84;
			2421: Pixel = 91;
			2422: Pixel = 97;
			2423: Pixel = 98;
			2424: Pixel = 100;
			2425: Pixel = 101;
			2426: Pixel = 103;
			2427: Pixel = 102;
			2428: Pixel = 103;
			2429: Pixel = 105;
			2430: Pixel = 107;
			2431: Pixel = 115;
			2432: Pixel = 117;
			2433: Pixel = 119;
			2434: Pixel = 120;
			2435: Pixel = 122;
			2436: Pixel = 123;
			2437: Pixel = 125;
			2438: Pixel = 125;
			2439: Pixel = 124;
			2440: Pixel = 125;
			2441: Pixel = 127;
			2442: Pixel = 128;
			2443: Pixel = 126;
			2444: Pixel = 126;
			2445: Pixel = 128;
			2446: Pixel = 128;
			2447: Pixel = 125;
			2448: Pixel = 120;
			2449: Pixel = 124;
			2450: Pixel = 130;
			2451: Pixel = 135;
			2452: Pixel = 134;
			2453: Pixel = 126;
			2454: Pixel = 132;
			2455: Pixel = 146;
			2456: Pixel = 142;
			2457: Pixel = 148;
			2458: Pixel = 145;
			2459: Pixel = 143;
			2460: Pixel = 148;
			2461: Pixel = 149;
			2462: Pixel = 154;
			2463: Pixel = 158;
			2464: Pixel = 162;
			2465: Pixel = 166;
			2466: Pixel = 174;
			2467: Pixel = 179;
			2468: Pixel = 175;
			2469: Pixel = 174;
			2470: Pixel = 176;
			2471: Pixel = 179;
			2472: Pixel = 180;
			2473: Pixel = 186;
			2474: Pixel = 192;
			2475: Pixel = 199;
			2476: Pixel = 194;
			2477: Pixel = 156;
			2478: Pixel = 116;
			2479: Pixel = 111;
			2480: Pixel = 122;
			2481: Pixel = 125;
			2482: Pixel = 127;
			2483: Pixel = 128;
			2484: Pixel = 124;
			2485: Pixel = 124;
			2486: Pixel = 126;
			2487: Pixel = 122;
			2488: Pixel = 122;
			2489: Pixel = 121;
			2490: Pixel = 118;
			2491: Pixel = 115;
			2492: Pixel = 113;
			2493: Pixel = 113;
			2494: Pixel = 111;
			2495: Pixel = 107;
			2496: Pixel = 110;
			2497: Pixel = 120;
			2498: Pixel = 133;
			2499: Pixel = 142;
			2500: Pixel = 145;
			2501: Pixel = 145;
			2502: Pixel = 144;
			2503: Pixel = 146;
			2504: Pixel = 148;
			2505: Pixel = 150;
			2506: Pixel = 152;
			2507: Pixel = 152;
			2508: Pixel = 152;
			2509: Pixel = 148;
			2510: Pixel = 149;
			2511: Pixel = 148;
			2512: Pixel = 146;
			2513: Pixel = 146;
			2514: Pixel = 146;
			2515: Pixel = 144;
			2516: Pixel = 143;
			2517: Pixel = 144;
			2518: Pixel = 141;
			2519: Pixel = 139;
			2520: Pixel = 139;
			2521: Pixel = 139;
			2522: Pixel = 141;
			2523: Pixel = 141;
			2524: Pixel = 140;
			2525: Pixel = 136;
			2526: Pixel = 148;
			2527: Pixel = 200;
			2528: Pixel = 219;
			2529: Pixel = 223;
			2530: Pixel = 226;
			2531: Pixel = 225;
			2532: Pixel = 181;
			2533: Pixel = 99;
			2534: Pixel = 49;
			2535: Pixel = 41;
			2536: Pixel = 43;
			2537: Pixel = 46;
			2538: Pixel = 50;
			2539: Pixel = 53;
			2540: Pixel = 54;
			2541: Pixel = 53;
			2542: Pixel = 53;
			2543: Pixel = 50;
			2544: Pixel = 45;
			2545: Pixel = 53;
			2546: Pixel = 50;
			2547: Pixel = 45;
			2548: Pixel = 44;
			2549: Pixel = 47;
			2550: Pixel = 160;
			2551: Pixel = 165;
			2552: Pixel = 171;
			2553: Pixel = 167;
			2554: Pixel = 156;
			2555: Pixel = 143;
			2556: Pixel = 122;
			2557: Pixel = 112;
			2558: Pixel = 131;
			2559: Pixel = 152;
			2560: Pixel = 161;
			2561: Pixel = 166;
			2562: Pixel = 165;
			2563: Pixel = 163;
			2564: Pixel = 164;
			2565: Pixel = 160;
			2566: Pixel = 151;
			2567: Pixel = 132;
			2568: Pixel = 100;
			2569: Pixel = 79;
			2570: Pixel = 82;
			2571: Pixel = 92;
			2572: Pixel = 95;
			2573: Pixel = 98;
			2574: Pixel = 99;
			2575: Pixel = 99;
			2576: Pixel = 99;
			2577: Pixel = 99;
			2578: Pixel = 102;
			2579: Pixel = 106;
			2580: Pixel = 106;
			2581: Pixel = 111;
			2582: Pixel = 114;
			2583: Pixel = 117;
			2584: Pixel = 118;
			2585: Pixel = 121;
			2586: Pixel = 122;
			2587: Pixel = 121;
			2588: Pixel = 122;
			2589: Pixel = 122;
			2590: Pixel = 123;
			2591: Pixel = 124;
			2592: Pixel = 126;
			2593: Pixel = 126;
			2594: Pixel = 127;
			2595: Pixel = 126;
			2596: Pixel = 121;
			2597: Pixel = 127;
			2598: Pixel = 142;
			2599: Pixel = 144;
			2600: Pixel = 149;
			2601: Pixel = 140;
			2602: Pixel = 127;
			2603: Pixel = 119;
			2604: Pixel = 128;
			2605: Pixel = 136;
			2606: Pixel = 137;
			2607: Pixel = 135;
			2608: Pixel = 138;
			2609: Pixel = 147;
			2610: Pixel = 148;
			2611: Pixel = 149;
			2612: Pixel = 152;
			2613: Pixel = 155;
			2614: Pixel = 165;
			2615: Pixel = 166;
			2616: Pixel = 169;
			2617: Pixel = 168;
			2618: Pixel = 174;
			2619: Pixel = 177;
			2620: Pixel = 175;
			2621: Pixel = 184;
			2622: Pixel = 187;
			2623: Pixel = 187;
			2624: Pixel = 190;
			2625: Pixel = 193;
			2626: Pixel = 195;
			2627: Pixel = 201;
			2628: Pixel = 182;
			2629: Pixel = 128;
			2630: Pixel = 110;
			2631: Pixel = 119;
			2632: Pixel = 121;
			2633: Pixel = 123;
			2634: Pixel = 120;
			2635: Pixel = 122;
			2636: Pixel = 122;
			2637: Pixel = 121;
			2638: Pixel = 122;
			2639: Pixel = 117;
			2640: Pixel = 114;
			2641: Pixel = 114;
			2642: Pixel = 112;
			2643: Pixel = 110;
			2644: Pixel = 106;
			2645: Pixel = 103;
			2646: Pixel = 109;
			2647: Pixel = 118;
			2648: Pixel = 132;
			2649: Pixel = 142;
			2650: Pixel = 146;
			2651: Pixel = 146;
			2652: Pixel = 144;
			2653: Pixel = 145;
			2654: Pixel = 148;
			2655: Pixel = 147;
			2656: Pixel = 149;
			2657: Pixel = 152;
			2658: Pixel = 152;
			2659: Pixel = 150;
			2660: Pixel = 145;
			2661: Pixel = 145;
			2662: Pixel = 144;
			2663: Pixel = 144;
			2664: Pixel = 145;
			2665: Pixel = 145;
			2666: Pixel = 143;
			2667: Pixel = 142;
			2668: Pixel = 141;
			2669: Pixel = 140;
			2670: Pixel = 140;
			2671: Pixel = 140;
			2672: Pixel = 140;
			2673: Pixel = 141;
			2674: Pixel = 141;
			2675: Pixel = 141;
			2676: Pixel = 134;
			2677: Pixel = 170;
			2678: Pixel = 213;
			2679: Pixel = 220;
			2680: Pixel = 225;
			2681: Pixel = 229;
			2682: Pixel = 215;
			2683: Pixel = 73;
			2684: Pixel = 34;
			2685: Pixel = 43;
			2686: Pixel = 45;
			2687: Pixel = 45;
			2688: Pixel = 51;
			2689: Pixel = 54;
			2690: Pixel = 51;
			2691: Pixel = 53;
			2692: Pixel = 50;
			2693: Pixel = 47;
			2694: Pixel = 51;
			2695: Pixel = 53;
			2696: Pixel = 47;
			2697: Pixel = 49;
			2698: Pixel = 46;
			2699: Pixel = 49;
			2700: Pixel = 163;
			2701: Pixel = 170;
			2702: Pixel = 170;
			2703: Pixel = 160;
			2704: Pixel = 150;
			2705: Pixel = 130;
			2706: Pixel = 101;
			2707: Pixel = 102;
			2708: Pixel = 132;
			2709: Pixel = 151;
			2710: Pixel = 162;
			2711: Pixel = 167;
			2712: Pixel = 165;
			2713: Pixel = 164;
			2714: Pixel = 165;
			2715: Pixel = 162;
			2716: Pixel = 151;
			2717: Pixel = 132;
			2718: Pixel = 102;
			2719: Pixel = 79;
			2720: Pixel = 79;
			2721: Pixel = 86;
			2722: Pixel = 90;
			2723: Pixel = 97;
			2724: Pixel = 97;
			2725: Pixel = 97;
			2726: Pixel = 98;
			2727: Pixel = 100;
			2728: Pixel = 102;
			2729: Pixel = 103;
			2730: Pixel = 106;
			2731: Pixel = 109;
			2732: Pixel = 113;
			2733: Pixel = 117;
			2734: Pixel = 116;
			2735: Pixel = 120;
			2736: Pixel = 120;
			2737: Pixel = 120;
			2738: Pixel = 123;
			2739: Pixel = 123;
			2740: Pixel = 122;
			2741: Pixel = 125;
			2742: Pixel = 125;
			2743: Pixel = 125;
			2744: Pixel = 125;
			2745: Pixel = 121;
			2746: Pixel = 141;
			2747: Pixel = 130;
			2748: Pixel = 137;
			2749: Pixel = 136;
			2750: Pixel = 127;
			2751: Pixel = 123;
			2752: Pixel = 123;
			2753: Pixel = 122;
			2754: Pixel = 126;
			2755: Pixel = 135;
			2756: Pixel = 131;
			2757: Pixel = 126;
			2758: Pixel = 137;
			2759: Pixel = 136;
			2760: Pixel = 141;
			2761: Pixel = 151;
			2762: Pixel = 150;
			2763: Pixel = 158;
			2764: Pixel = 161;
			2765: Pixel = 160;
			2766: Pixel = 167;
			2767: Pixel = 170;
			2768: Pixel = 176;
			2769: Pixel = 181;
			2770: Pixel = 185;
			2771: Pixel = 184;
			2772: Pixel = 183;
			2773: Pixel = 187;
			2774: Pixel = 188;
			2775: Pixel = 190;
			2776: Pixel = 192;
			2777: Pixel = 195;
			2778: Pixel = 201;
			2779: Pixel = 197;
			2780: Pixel = 156;
			2781: Pixel = 111;
			2782: Pixel = 107;
			2783: Pixel = 117;
			2784: Pixel = 118;
			2785: Pixel = 120;
			2786: Pixel = 120;
			2787: Pixel = 119;
			2788: Pixel = 119;
			2789: Pixel = 118;
			2790: Pixel = 116;
			2791: Pixel = 113;
			2792: Pixel = 111;
			2793: Pixel = 108;
			2794: Pixel = 106;
			2795: Pixel = 101;
			2796: Pixel = 106;
			2797: Pixel = 118;
			2798: Pixel = 133;
			2799: Pixel = 141;
			2800: Pixel = 148;
			2801: Pixel = 147;
			2802: Pixel = 144;
			2803: Pixel = 144;
			2804: Pixel = 147;
			2805: Pixel = 146;
			2806: Pixel = 146;
			2807: Pixel = 149;
			2808: Pixel = 150;
			2809: Pixel = 153;
			2810: Pixel = 147;
			2811: Pixel = 142;
			2812: Pixel = 140;
			2813: Pixel = 142;
			2814: Pixel = 144;
			2815: Pixel = 145;
			2816: Pixel = 143;
			2817: Pixel = 142;
			2818: Pixel = 144;
			2819: Pixel = 141;
			2820: Pixel = 140;
			2821: Pixel = 141;
			2822: Pixel = 140;
			2823: Pixel = 143;
			2824: Pixel = 144;
			2825: Pixel = 142;
			2826: Pixel = 138;
			2827: Pixel = 143;
			2828: Pixel = 192;
			2829: Pixel = 219;
			2830: Pixel = 224;
			2831: Pixel = 236;
			2832: Pixel = 169;
			2833: Pixel = 39;
			2834: Pixel = 39;
			2835: Pixel = 44;
			2836: Pixel = 46;
			2837: Pixel = 50;
			2838: Pixel = 53;
			2839: Pixel = 52;
			2840: Pixel = 54;
			2841: Pixel = 49;
			2842: Pixel = 43;
			2843: Pixel = 46;
			2844: Pixel = 54;
			2845: Pixel = 48;
			2846: Pixel = 43;
			2847: Pixel = 46;
			2848: Pixel = 50;
			2849: Pixel = 54;
			2850: Pixel = 169;
			2851: Pixel = 174;
			2852: Pixel = 166;
			2853: Pixel = 155;
			2854: Pixel = 142;
			2855: Pixel = 113;
			2856: Pixel = 81;
			2857: Pixel = 99;
			2858: Pixel = 134;
			2859: Pixel = 152;
			2860: Pixel = 164;
			2861: Pixel = 166;
			2862: Pixel = 165;
			2863: Pixel = 164;
			2864: Pixel = 163;
			2865: Pixel = 160;
			2866: Pixel = 148;
			2867: Pixel = 131;
			2868: Pixel = 101;
			2869: Pixel = 75;
			2870: Pixel = 77;
			2871: Pixel = 85;
			2872: Pixel = 92;
			2873: Pixel = 94;
			2874: Pixel = 94;
			2875: Pixel = 97;
			2876: Pixel = 99;
			2877: Pixel = 99;
			2878: Pixel = 101;
			2879: Pixel = 103;
			2880: Pixel = 104;
			2881: Pixel = 105;
			2882: Pixel = 109;
			2883: Pixel = 115;
			2884: Pixel = 115;
			2885: Pixel = 117;
			2886: Pixel = 115;
			2887: Pixel = 121;
			2888: Pixel = 124;
			2889: Pixel = 123;
			2890: Pixel = 123;
			2891: Pixel = 123;
			2892: Pixel = 124;
			2893: Pixel = 124;
			2894: Pixel = 118;
			2895: Pixel = 135;
			2896: Pixel = 150;
			2897: Pixel = 101;
			2898: Pixel = 120;
			2899: Pixel = 120;
			2900: Pixel = 119;
			2901: Pixel = 122;
			2902: Pixel = 122;
			2903: Pixel = 120;
			2904: Pixel = 128;
			2905: Pixel = 133;
			2906: Pixel = 129;
			2907: Pixel = 128;
			2908: Pixel = 134;
			2909: Pixel = 136;
			2910: Pixel = 138;
			2911: Pixel = 142;
			2912: Pixel = 145;
			2913: Pixel = 153;
			2914: Pixel = 153;
			2915: Pixel = 161;
			2916: Pixel = 172;
			2917: Pixel = 172;
			2918: Pixel = 175;
			2919: Pixel = 184;
			2920: Pixel = 184;
			2921: Pixel = 185;
			2922: Pixel = 184;
			2923: Pixel = 189;
			2924: Pixel = 186;
			2925: Pixel = 187;
			2926: Pixel = 193;
			2927: Pixel = 195;
			2928: Pixel = 194;
			2929: Pixel = 196;
			2930: Pixel = 198;
			2931: Pixel = 177;
			2932: Pixel = 124;
			2933: Pixel = 100;
			2934: Pixel = 111;
			2935: Pixel = 116;
			2936: Pixel = 114;
			2937: Pixel = 116;
			2938: Pixel = 117;
			2939: Pixel = 116;
			2940: Pixel = 115;
			2941: Pixel = 111;
			2942: Pixel = 110;
			2943: Pixel = 108;
			2944: Pixel = 106;
			2945: Pixel = 102;
			2946: Pixel = 105;
			2947: Pixel = 118;
			2948: Pixel = 134;
			2949: Pixel = 144;
			2950: Pixel = 149;
			2951: Pixel = 150;
			2952: Pixel = 146;
			2953: Pixel = 144;
			2954: Pixel = 144;
			2955: Pixel = 144;
			2956: Pixel = 143;
			2957: Pixel = 142;
			2958: Pixel = 146;
			2959: Pixel = 150;
			2960: Pixel = 148;
			2961: Pixel = 141;
			2962: Pixel = 140;
			2963: Pixel = 141;
			2964: Pixel = 142;
			2965: Pixel = 145;
			2966: Pixel = 143;
			2967: Pixel = 142;
			2968: Pixel = 142;
			2969: Pixel = 141;
			2970: Pixel = 140;
			2971: Pixel = 141;
			2972: Pixel = 140;
			2973: Pixel = 144;
			2974: Pixel = 143;
			2975: Pixel = 143;
			2976: Pixel = 143;
			2977: Pixel = 140;
			2978: Pixel = 159;
			2979: Pixel = 212;
			2980: Pixel = 231;
			2981: Pixel = 195;
			2982: Pixel = 65;
			2983: Pixel = 34;
			2984: Pixel = 43;
			2985: Pixel = 43;
			2986: Pixel = 48;
			2987: Pixel = 54;
			2988: Pixel = 54;
			2989: Pixel = 55;
			2990: Pixel = 53;
			2991: Pixel = 43;
			2992: Pixel = 45;
			2993: Pixel = 51;
			2994: Pixel = 48;
			2995: Pixel = 44;
			2996: Pixel = 45;
			2997: Pixel = 52;
			2998: Pixel = 53;
			2999: Pixel = 37;
			3000: Pixel = 172;
			3001: Pixel = 171;
			3002: Pixel = 160;
			3003: Pixel = 149;
			3004: Pixel = 127;
			3005: Pixel = 90;
			3006: Pixel = 74;
			3007: Pixel = 102;
			3008: Pixel = 131;
			3009: Pixel = 149;
			3010: Pixel = 163;
			3011: Pixel = 167;
			3012: Pixel = 164;
			3013: Pixel = 164;
			3014: Pixel = 164;
			3015: Pixel = 159;
			3016: Pixel = 145;
			3017: Pixel = 130;
			3018: Pixel = 100;
			3019: Pixel = 75;
			3020: Pixel = 77;
			3021: Pixel = 87;
			3022: Pixel = 91;
			3023: Pixel = 97;
			3024: Pixel = 101;
			3025: Pixel = 100;
			3026: Pixel = 100;
			3027: Pixel = 99;
			3028: Pixel = 101;
			3029: Pixel = 101;
			3030: Pixel = 104;
			3031: Pixel = 108;
			3032: Pixel = 111;
			3033: Pixel = 115;
			3034: Pixel = 112;
			3035: Pixel = 115;
			3036: Pixel = 117;
			3037: Pixel = 119;
			3038: Pixel = 119;
			3039: Pixel = 120;
			3040: Pixel = 123;
			3041: Pixel = 124;
			3042: Pixel = 124;
			3043: Pixel = 123;
			3044: Pixel = 122;
			3045: Pixel = 131;
			3046: Pixel = 115;
			3047: Pixel = 109;
			3048: Pixel = 120;
			3049: Pixel = 120;
			3050: Pixel = 119;
			3051: Pixel = 124;
			3052: Pixel = 121;
			3053: Pixel = 121;
			3054: Pixel = 129;
			3055: Pixel = 133;
			3056: Pixel = 129;
			3057: Pixel = 129;
			3058: Pixel = 136;
			3059: Pixel = 134;
			3060: Pixel = 131;
			3061: Pixel = 137;
			3062: Pixel = 138;
			3063: Pixel = 147;
			3064: Pixel = 156;
			3065: Pixel = 164;
			3066: Pixel = 173;
			3067: Pixel = 176;
			3068: Pixel = 175;
			3069: Pixel = 178;
			3070: Pixel = 180;
			3071: Pixel = 182;
			3072: Pixel = 184;
			3073: Pixel = 188;
			3074: Pixel = 191;
			3075: Pixel = 190;
			3076: Pixel = 192;
			3077: Pixel = 196;
			3078: Pixel = 197;
			3079: Pixel = 195;
			3080: Pixel = 193;
			3081: Pixel = 204;
			3082: Pixel = 200;
			3083: Pixel = 141;
			3084: Pixel = 96;
			3085: Pixel = 101;
			3086: Pixel = 107;
			3087: Pixel = 110;
			3088: Pixel = 113;
			3089: Pixel = 113;
			3090: Pixel = 113;
			3091: Pixel = 110;
			3092: Pixel = 109;
			3093: Pixel = 107;
			3094: Pixel = 107;
			3095: Pixel = 101;
			3096: Pixel = 104;
			3097: Pixel = 117;
			3098: Pixel = 134;
			3099: Pixel = 145;
			3100: Pixel = 151;
			3101: Pixel = 151;
			3102: Pixel = 149;
			3103: Pixel = 148;
			3104: Pixel = 144;
			3105: Pixel = 140;
			3106: Pixel = 140;
			3107: Pixel = 138;
			3108: Pixel = 138;
			3109: Pixel = 145;
			3110: Pixel = 149;
			3111: Pixel = 144;
			3112: Pixel = 142;
			3113: Pixel = 142;
			3114: Pixel = 144;
			3115: Pixel = 145;
			3116: Pixel = 144;
			3117: Pixel = 142;
			3118: Pixel = 142;
			3119: Pixel = 142;
			3120: Pixel = 141;
			3121: Pixel = 143;
			3122: Pixel = 143;
			3123: Pixel = 144;
			3124: Pixel = 144;
			3125: Pixel = 145;
			3126: Pixel = 146;
			3127: Pixel = 149;
			3128: Pixel = 148;
			3129: Pixel = 194;
			3130: Pixel = 184;
			3131: Pixel = 73;
			3132: Pixel = 37;
			3133: Pixel = 46;
			3134: Pixel = 44;
			3135: Pixel = 45;
			3136: Pixel = 49;
			3137: Pixel = 50;
			3138: Pixel = 53;
			3139: Pixel = 54;
			3140: Pixel = 47;
			3141: Pixel = 50;
			3142: Pixel = 53;
			3143: Pixel = 52;
			3144: Pixel = 45;
			3145: Pixel = 45;
			3146: Pixel = 55;
			3147: Pixel = 65;
			3148: Pixel = 39;
			3149: Pixel = 26;
			3150: Pixel = 172;
			3151: Pixel = 166;
			3152: Pixel = 155;
			3153: Pixel = 139;
			3154: Pixel = 108;
			3155: Pixel = 76;
			3156: Pixel = 79;
			3157: Pixel = 104;
			3158: Pixel = 131;
			3159: Pixel = 150;
			3160: Pixel = 163;
			3161: Pixel = 168;
			3162: Pixel = 166;
			3163: Pixel = 164;
			3164: Pixel = 163;
			3165: Pixel = 158;
			3166: Pixel = 146;
			3167: Pixel = 130;
			3168: Pixel = 98;
			3169: Pixel = 72;
			3170: Pixel = 77;
			3171: Pixel = 87;
			3172: Pixel = 92;
			3173: Pixel = 98;
			3174: Pixel = 99;
			3175: Pixel = 102;
			3176: Pixel = 100;
			3177: Pixel = 98;
			3178: Pixel = 100;
			3179: Pixel = 99;
			3180: Pixel = 104;
			3181: Pixel = 108;
			3182: Pixel = 110;
			3183: Pixel = 113;
			3184: Pixel = 115;
			3185: Pixel = 115;
			3186: Pixel = 116;
			3187: Pixel = 119;
			3188: Pixel = 119;
			3189: Pixel = 120;
			3190: Pixel = 121;
			3191: Pixel = 123;
			3192: Pixel = 124;
			3193: Pixel = 118;
			3194: Pixel = 141;
			3195: Pixel = 129;
			3196: Pixel = 109;
			3197: Pixel = 117;
			3198: Pixel = 113;
			3199: Pixel = 110;
			3200: Pixel = 117;
			3201: Pixel = 121;
			3202: Pixel = 126;
			3203: Pixel = 124;
			3204: Pixel = 130;
			3205: Pixel = 127;
			3206: Pixel = 133;
			3207: Pixel = 135;
			3208: Pixel = 137;
			3209: Pixel = 130;
			3210: Pixel = 135;
			3211: Pixel = 139;
			3212: Pixel = 140;
			3213: Pixel = 145;
			3214: Pixel = 150;
			3215: Pixel = 159;
			3216: Pixel = 164;
			3217: Pixel = 167;
			3218: Pixel = 172;
			3219: Pixel = 180;
			3220: Pixel = 182;
			3221: Pixel = 183;
			3222: Pixel = 189;
			3223: Pixel = 191;
			3224: Pixel = 191;
			3225: Pixel = 192;
			3226: Pixel = 194;
			3227: Pixel = 196;
			3228: Pixel = 195;
			3229: Pixel = 195;
			3230: Pixel = 198;
			3231: Pixel = 197;
			3232: Pixel = 198;
			3233: Pixel = 203;
			3234: Pixel = 148;
			3235: Pixel = 97;
			3236: Pixel = 92;
			3237: Pixel = 98;
			3238: Pixel = 107;
			3239: Pixel = 111;
			3240: Pixel = 110;
			3241: Pixel = 108;
			3242: Pixel = 106;
			3243: Pixel = 108;
			3244: Pixel = 107;
			3245: Pixel = 101;
			3246: Pixel = 102;
			3247: Pixel = 115;
			3248: Pixel = 135;
			3249: Pixel = 148;
			3250: Pixel = 152;
			3251: Pixel = 154;
			3252: Pixel = 153;
			3253: Pixel = 150;
			3254: Pixel = 146;
			3255: Pixel = 137;
			3256: Pixel = 132;
			3257: Pixel = 130;
			3258: Pixel = 130;
			3259: Pixel = 138;
			3260: Pixel = 148;
			3261: Pixel = 148;
			3262: Pixel = 143;
			3263: Pixel = 142;
			3264: Pixel = 145;
			3265: Pixel = 147;
			3266: Pixel = 143;
			3267: Pixel = 142;
			3268: Pixel = 142;
			3269: Pixel = 141;
			3270: Pixel = 143;
			3271: Pixel = 145;
			3272: Pixel = 144;
			3273: Pixel = 145;
			3274: Pixel = 146;
			3275: Pixel = 148;
			3276: Pixel = 148;
			3277: Pixel = 149;
			3278: Pixel = 158;
			3279: Pixel = 145;
			3280: Pixel = 67;
			3281: Pixel = 38;
			3282: Pixel = 47;
			3283: Pixel = 42;
			3284: Pixel = 46;
			3285: Pixel = 52;
			3286: Pixel = 52;
			3287: Pixel = 51;
			3288: Pixel = 51;
			3289: Pixel = 44;
			3290: Pixel = 44;
			3291: Pixel = 58;
			3292: Pixel = 53;
			3293: Pixel = 47;
			3294: Pixel = 48;
			3295: Pixel = 55;
			3296: Pixel = 68;
			3297: Pixel = 51;
			3298: Pixel = 28;
			3299: Pixel = 77;
			3300: Pixel = 168;
			3301: Pixel = 161;
			3302: Pixel = 149;
			3303: Pixel = 122;
			3304: Pixel = 88;
			3305: Pixel = 81;
			3306: Pixel = 80;
			3307: Pixel = 105;
			3308: Pixel = 131;
			3309: Pixel = 150;
			3310: Pixel = 164;
			3311: Pixel = 167;
			3312: Pixel = 168;
			3313: Pixel = 165;
			3314: Pixel = 163;
			3315: Pixel = 158;
			3316: Pixel = 148;
			3317: Pixel = 129;
			3318: Pixel = 98;
			3319: Pixel = 74;
			3320: Pixel = 79;
			3321: Pixel = 86;
			3322: Pixel = 93;
			3323: Pixel = 100;
			3324: Pixel = 98;
			3325: Pixel = 99;
			3326: Pixel = 99;
			3327: Pixel = 100;
			3328: Pixel = 100;
			3329: Pixel = 101;
			3330: Pixel = 103;
			3331: Pixel = 106;
			3332: Pixel = 110;
			3333: Pixel = 113;
			3334: Pixel = 116;
			3335: Pixel = 113;
			3336: Pixel = 116;
			3337: Pixel = 120;
			3338: Pixel = 118;
			3339: Pixel = 119;
			3340: Pixel = 122;
			3341: Pixel = 121;
			3342: Pixel = 123;
			3343: Pixel = 124;
			3344: Pixel = 151;
			3345: Pixel = 118;
			3346: Pixel = 111;
			3347: Pixel = 108;
			3348: Pixel = 107;
			3349: Pixel = 115;
			3350: Pixel = 118;
			3351: Pixel = 118;
			3352: Pixel = 123;
			3353: Pixel = 126;
			3354: Pixel = 124;
			3355: Pixel = 129;
			3356: Pixel = 131;
			3357: Pixel = 131;
			3358: Pixel = 137;
			3359: Pixel = 138;
			3360: Pixel = 136;
			3361: Pixel = 137;
			3362: Pixel = 136;
			3363: Pixel = 147;
			3364: Pixel = 147;
			3365: Pixel = 152;
			3366: Pixel = 159;
			3367: Pixel = 168;
			3368: Pixel = 177;
			3369: Pixel = 181;
			3370: Pixel = 184;
			3371: Pixel = 186;
			3372: Pixel = 186;
			3373: Pixel = 189;
			3374: Pixel = 190;
			3375: Pixel = 191;
			3376: Pixel = 196;
			3377: Pixel = 196;
			3378: Pixel = 194;
			3379: Pixel = 189;
			3380: Pixel = 189;
			3381: Pixel = 190;
			3382: Pixel = 195;
			3383: Pixel = 208;
			3384: Pixel = 218;
			3385: Pixel = 209;
			3386: Pixel = 166;
			3387: Pixel = 89;
			3388: Pixel = 97;
			3389: Pixel = 107;
			3390: Pixel = 107;
			3391: Pixel = 105;
			3392: Pixel = 103;
			3393: Pixel = 105;
			3394: Pixel = 104;
			3395: Pixel = 99;
			3396: Pixel = 103;
			3397: Pixel = 116;
			3398: Pixel = 137;
			3399: Pixel = 149;
			3400: Pixel = 154;
			3401: Pixel = 156;
			3402: Pixel = 155;
			3403: Pixel = 152;
			3404: Pixel = 149;
			3405: Pixel = 137;
			3406: Pixel = 124;
			3407: Pixel = 116;
			3408: Pixel = 118;
			3409: Pixel = 131;
			3410: Pixel = 143;
			3411: Pixel = 149;
			3412: Pixel = 145;
			3413: Pixel = 144;
			3414: Pixel = 146;
			3415: Pixel = 148;
			3416: Pixel = 144;
			3417: Pixel = 142;
			3418: Pixel = 142;
			3419: Pixel = 142;
			3420: Pixel = 144;
			3421: Pixel = 144;
			3422: Pixel = 144;
			3423: Pixel = 146;
			3424: Pixel = 145;
			3425: Pixel = 148;
			3426: Pixel = 149;
			3427: Pixel = 155;
			3428: Pixel = 154;
			3429: Pixel = 81;
			3430: Pixel = 39;
			3431: Pixel = 46;
			3432: Pixel = 43;
			3433: Pixel = 42;
			3434: Pixel = 48;
			3435: Pixel = 53;
			3436: Pixel = 54;
			3437: Pixel = 49;
			3438: Pixel = 44;
			3439: Pixel = 45;
			3440: Pixel = 54;
			3441: Pixel = 54;
			3442: Pixel = 49;
			3443: Pixel = 48;
			3444: Pixel = 52;
			3445: Pixel = 69;
			3446: Pixel = 55;
			3447: Pixel = 30;
			3448: Pixel = 67;
			3449: Pixel = 150;
			3450: Pixel = 162;
			3451: Pixel = 153;
			3452: Pixel = 135;
			3453: Pixel = 103;
			3454: Pixel = 80;
			3455: Pixel = 85;
			3456: Pixel = 82;
			3457: Pixel = 105;
			3458: Pixel = 133;
			3459: Pixel = 150;
			3460: Pixel = 162;
			3461: Pixel = 167;
			3462: Pixel = 167;
			3463: Pixel = 167;
			3464: Pixel = 163;
			3465: Pixel = 159;
			3466: Pixel = 148;
			3467: Pixel = 128;
			3468: Pixel = 98;
			3469: Pixel = 75;
			3470: Pixel = 77;
			3471: Pixel = 87;
			3472: Pixel = 93;
			3473: Pixel = 99;
			3474: Pixel = 98;
			3475: Pixel = 99;
			3476: Pixel = 100;
			3477: Pixel = 99;
			3478: Pixel = 101;
			3479: Pixel = 102;
			3480: Pixel = 104;
			3481: Pixel = 108;
			3482: Pixel = 111;
			3483: Pixel = 114;
			3484: Pixel = 115;
			3485: Pixel = 114;
			3486: Pixel = 117;
			3487: Pixel = 120;
			3488: Pixel = 121;
			3489: Pixel = 122;
			3490: Pixel = 121;
			3491: Pixel = 120;
			3492: Pixel = 122;
			3493: Pixel = 131;
			3494: Pixel = 126;
			3495: Pixel = 109;
			3496: Pixel = 108;
			3497: Pixel = 108;
			3498: Pixel = 113;
			3499: Pixel = 120;
			3500: Pixel = 115;
			3501: Pixel = 118;
			3502: Pixel = 124;
			3503: Pixel = 123;
			3504: Pixel = 123;
			3505: Pixel = 129;
			3506: Pixel = 125;
			3507: Pixel = 127;
			3508: Pixel = 133;
			3509: Pixel = 133;
			3510: Pixel = 134;
			3511: Pixel = 133;
			3512: Pixel = 141;
			3513: Pixel = 144;
			3514: Pixel = 146;
			3515: Pixel = 155;
			3516: Pixel = 160;
			3517: Pixel = 172;
			3518: Pixel = 180;
			3519: Pixel = 185;
			3520: Pixel = 186;
			3521: Pixel = 183;
			3522: Pixel = 185;
			3523: Pixel = 187;
			3524: Pixel = 192;
			3525: Pixel = 193;
			3526: Pixel = 190;
			3527: Pixel = 186;
			3528: Pixel = 186;
			3529: Pixel = 192;
			3530: Pixel = 202;
			3531: Pixel = 209;
			3532: Pixel = 215;
			3533: Pixel = 214;
			3534: Pixel = 217;
			3535: Pixel = 228;
			3536: Pixel = 237;
			3537: Pixel = 141;
			3538: Pixel = 74;
			3539: Pixel = 99;
			3540: Pixel = 103;
			3541: Pixel = 102;
			3542: Pixel = 101;
			3543: Pixel = 102;
			3544: Pixel = 102;
			3545: Pixel = 98;
			3546: Pixel = 103;
			3547: Pixel = 115;
			3548: Pixel = 135;
			3549: Pixel = 146;
			3550: Pixel = 153;
			3551: Pixel = 155;
			3552: Pixel = 154;
			3553: Pixel = 153;
			3554: Pixel = 152;
			3555: Pixel = 140;
			3556: Pixel = 120;
			3557: Pixel = 100;
			3558: Pixel = 98;
			3559: Pixel = 115;
			3560: Pixel = 134;
			3561: Pixel = 146;
			3562: Pixel = 149;
			3563: Pixel = 144;
			3564: Pixel = 143;
			3565: Pixel = 145;
			3566: Pixel = 145;
			3567: Pixel = 142;
			3568: Pixel = 143;
			3569: Pixel = 144;
			3570: Pixel = 144;
			3571: Pixel = 143;
			3572: Pixel = 143;
			3573: Pixel = 145;
			3574: Pixel = 147;
			3575: Pixel = 148;
			3576: Pixel = 152;
			3577: Pixel = 158;
			3578: Pixel = 102;
			3579: Pixel = 45;
			3580: Pixel = 46;
			3581: Pixel = 43;
			3582: Pixel = 45;
			3583: Pixel = 47;
			3584: Pixel = 52;
			3585: Pixel = 51;
			3586: Pixel = 51;
			3587: Pixel = 46;
			3588: Pixel = 43;
			3589: Pixel = 55;
			3590: Pixel = 55;
			3591: Pixel = 47;
			3592: Pixel = 46;
			3593: Pixel = 48;
			3594: Pixel = 66;
			3595: Pixel = 79;
			3596: Pixel = 42;
			3597: Pixel = 60;
			3598: Pixel = 131;
			3599: Pixel = 165;
			3600: Pixel = 157;
			3601: Pixel = 145;
			3602: Pixel = 117;
			3603: Pixel = 86;
			3604: Pixel = 82;
			3605: Pixel = 85;
			3606: Pixel = 85;
			3607: Pixel = 105;
			3608: Pixel = 132;
			3609: Pixel = 150;
			3610: Pixel = 161;
			3611: Pixel = 167;
			3612: Pixel = 167;
			3613: Pixel = 167;
			3614: Pixel = 164;
			3615: Pixel = 157;
			3616: Pixel = 145;
			3617: Pixel = 125;
			3618: Pixel = 98;
			3619: Pixel = 76;
			3620: Pixel = 78;
			3621: Pixel = 89;
			3622: Pixel = 94;
			3623: Pixel = 96;
			3624: Pixel = 101;
			3625: Pixel = 98;
			3626: Pixel = 100;
			3627: Pixel = 101;
			3628: Pixel = 99;
			3629: Pixel = 102;
			3630: Pixel = 103;
			3631: Pixel = 108;
			3632: Pixel = 112;
			3633: Pixel = 113;
			3634: Pixel = 114;
			3635: Pixel = 116;
			3636: Pixel = 118;
			3637: Pixel = 121;
			3638: Pixel = 121;
			3639: Pixel = 121;
			3640: Pixel = 121;
			3641: Pixel = 122;
			3642: Pixel = 126;
			3643: Pixel = 126;
			3644: Pixel = 109;
			3645: Pixel = 108;
			3646: Pixel = 110;
			3647: Pixel = 115;
			3648: Pixel = 119;
			3649: Pixel = 118;
			3650: Pixel = 119;
			3651: Pixel = 121;
			3652: Pixel = 121;
			3653: Pixel = 119;
			3654: Pixel = 120;
			3655: Pixel = 121;
			3656: Pixel = 127;
			3657: Pixel = 131;
			3658: Pixel = 135;
			3659: Pixel = 133;
			3660: Pixel = 134;
			3661: Pixel = 132;
			3662: Pixel = 139;
			3663: Pixel = 136;
			3664: Pixel = 142;
			3665: Pixel = 152;
			3666: Pixel = 160;
			3667: Pixel = 168;
			3668: Pixel = 182;
			3669: Pixel = 183;
			3670: Pixel = 185;
			3671: Pixel = 187;
			3672: Pixel = 190;
			3673: Pixel = 187;
			3674: Pixel = 184;
			3675: Pixel = 177;
			3676: Pixel = 179;
			3677: Pixel = 194;
			3678: Pixel = 206;
			3679: Pixel = 213;
			3680: Pixel = 211;
			3681: Pixel = 210;
			3682: Pixel = 210;
			3683: Pixel = 209;
			3684: Pixel = 209;
			3685: Pixel = 215;
			3686: Pixel = 226;
			3687: Pixel = 214;
			3688: Pixel = 103;
			3689: Pixel = 80;
			3690: Pixel = 98;
			3691: Pixel = 99;
			3692: Pixel = 100;
			3693: Pixel = 99;
			3694: Pixel = 100;
			3695: Pixel = 95;
			3696: Pixel = 99;
			3697: Pixel = 115;
			3698: Pixel = 133;
			3699: Pixel = 145;
			3700: Pixel = 153;
			3701: Pixel = 154;
			3702: Pixel = 152;
			3703: Pixel = 153;
			3704: Pixel = 151;
			3705: Pixel = 142;
			3706: Pixel = 124;
			3707: Pixel = 90;
			3708: Pixel = 73;
			3709: Pixel = 91;
			3710: Pixel = 124;
			3711: Pixel = 139;
			3712: Pixel = 147;
			3713: Pixel = 146;
			3714: Pixel = 143;
			3715: Pixel = 147;
			3716: Pixel = 145;
			3717: Pixel = 142;
			3718: Pixel = 144;
			3719: Pixel = 142;
			3720: Pixel = 144;
			3721: Pixel = 145;
			3722: Pixel = 144;
			3723: Pixel = 146;
			3724: Pixel = 147;
			3725: Pixel = 148;
			3726: Pixel = 159;
			3727: Pixel = 126;
			3728: Pixel = 50;
			3729: Pixel = 39;
			3730: Pixel = 40;
			3731: Pixel = 43;
			3732: Pixel = 47;
			3733: Pixel = 52;
			3734: Pixel = 53;
			3735: Pixel = 52;
			3736: Pixel = 48;
			3737: Pixel = 43;
			3738: Pixel = 48;
			3739: Pixel = 56;
			3740: Pixel = 47;
			3741: Pixel = 47;
			3742: Pixel = 48;
			3743: Pixel = 59;
			3744: Pixel = 74;
			3745: Pixel = 63;
			3746: Pixel = 63;
			3747: Pixel = 122;
			3748: Pixel = 153;
			3749: Pixel = 158;
			3750: Pixel = 148;
			3751: Pixel = 129;
			3752: Pixel = 94;
			3753: Pixel = 81;
			3754: Pixel = 89;
			3755: Pixel = 88;
			3756: Pixel = 85;
			3757: Pixel = 105;
			3758: Pixel = 132;
			3759: Pixel = 150;
			3760: Pixel = 162;
			3761: Pixel = 168;
			3762: Pixel = 167;
			3763: Pixel = 166;
			3764: Pixel = 165;
			3765: Pixel = 157;
			3766: Pixel = 144;
			3767: Pixel = 126;
			3768: Pixel = 101;
			3769: Pixel = 79;
			3770: Pixel = 79;
			3771: Pixel = 88;
			3772: Pixel = 93;
			3773: Pixel = 96;
			3774: Pixel = 98;
			3775: Pixel = 99;
			3776: Pixel = 101;
			3777: Pixel = 105;
			3778: Pixel = 101;
			3779: Pixel = 100;
			3780: Pixel = 103;
			3781: Pixel = 108;
			3782: Pixel = 110;
			3783: Pixel = 114;
			3784: Pixel = 115;
			3785: Pixel = 116;
			3786: Pixel = 117;
			3787: Pixel = 119;
			3788: Pixel = 120;
			3789: Pixel = 121;
			3790: Pixel = 123;
			3791: Pixel = 125;
			3792: Pixel = 126;
			3793: Pixel = 113;
			3794: Pixel = 104;
			3795: Pixel = 108;
			3796: Pixel = 113;
			3797: Pixel = 115;
			3798: Pixel = 116;
			3799: Pixel = 121;
			3800: Pixel = 120;
			3801: Pixel = 121;
			3802: Pixel = 119;
			3803: Pixel = 116;
			3804: Pixel = 119;
			3805: Pixel = 128;
			3806: Pixel = 130;
			3807: Pixel = 133;
			3808: Pixel = 139;
			3809: Pixel = 136;
			3810: Pixel = 135;
			3811: Pixel = 136;
			3812: Pixel = 140;
			3813: Pixel = 139;
			3814: Pixel = 145;
			3815: Pixel = 154;
			3816: Pixel = 158;
			3817: Pixel = 168;
			3818: Pixel = 177;
			3819: Pixel = 180;
			3820: Pixel = 181;
			3821: Pixel = 189;
			3822: Pixel = 185;
			3823: Pixel = 167;
			3824: Pixel = 174;
			3825: Pixel = 195;
			3826: Pixel = 210;
			3827: Pixel = 213;
			3828: Pixel = 205;
			3829: Pixel = 205;
			3830: Pixel = 207;
			3831: Pixel = 207;
			3832: Pixel = 205;
			3833: Pixel = 210;
			3834: Pixel = 207;
			3835: Pixel = 209;
			3836: Pixel = 216;
			3837: Pixel = 229;
			3838: Pixel = 190;
			3839: Pixel = 85;
			3840: Pixel = 82;
			3841: Pixel = 93;
			3842: Pixel = 97;
			3843: Pixel = 98;
			3844: Pixel = 97;
			3845: Pixel = 94;
			3846: Pixel = 98;
			3847: Pixel = 114;
			3848: Pixel = 131;
			3849: Pixel = 146;
			3850: Pixel = 155;
			3851: Pixel = 153;
			3852: Pixel = 152;
			3853: Pixel = 153;
			3854: Pixel = 150;
			3855: Pixel = 142;
			3856: Pixel = 127;
			3857: Pixel = 89;
			3858: Pixel = 53;
			3859: Pixel = 68;
			3860: Pixel = 109;
			3861: Pixel = 131;
			3862: Pixel = 144;
			3863: Pixel = 149;
			3864: Pixel = 145;
			3865: Pixel = 144;
			3866: Pixel = 146;
			3867: Pixel = 142;
			3868: Pixel = 144;
			3869: Pixel = 143;
			3870: Pixel = 144;
			3871: Pixel = 144;
			3872: Pixel = 142;
			3873: Pixel = 144;
			3874: Pixel = 147;
			3875: Pixel = 155;
			3876: Pixel = 147;
			3877: Pixel = 66;
			3878: Pixel = 35;
			3879: Pixel = 42;
			3880: Pixel = 41;
			3881: Pixel = 47;
			3882: Pixel = 55;
			3883: Pixel = 54;
			3884: Pixel = 53;
			3885: Pixel = 52;
			3886: Pixel = 41;
			3887: Pixel = 49;
			3888: Pixel = 56;
			3889: Pixel = 47;
			3890: Pixel = 43;
			3891: Pixel = 54;
			3892: Pixel = 65;
			3893: Pixel = 71;
			3894: Pixel = 72;
			3895: Pixel = 71;
			3896: Pixel = 119;
			3897: Pixel = 150;
			3898: Pixel = 146;
			3899: Pixel = 146;
			3900: Pixel = 137;
			3901: Pixel = 108;
			3902: Pixel = 82;
			3903: Pixel = 87;
			3904: Pixel = 90;
			3905: Pixel = 87;
			3906: Pixel = 85;
			3907: Pixel = 104;
			3908: Pixel = 131;
			3909: Pixel = 149;
			3910: Pixel = 160;
			3911: Pixel = 166;
			3912: Pixel = 166;
			3913: Pixel = 165;
			3914: Pixel = 165;
			3915: Pixel = 157;
			3916: Pixel = 144;
			3917: Pixel = 126;
			3918: Pixel = 99;
			3919: Pixel = 76;
			3920: Pixel = 79;
			3921: Pixel = 89;
			3922: Pixel = 94;
			3923: Pixel = 96;
			3924: Pixel = 97;
			3925: Pixel = 101;
			3926: Pixel = 101;
			3927: Pixel = 102;
			3928: Pixel = 99;
			3929: Pixel = 100;
			3930: Pixel = 105;
			3931: Pixel = 108;
			3932: Pixel = 108;
			3933: Pixel = 113;
			3934: Pixel = 116;
			3935: Pixel = 115;
			3936: Pixel = 119;
			3937: Pixel = 122;
			3938: Pixel = 121;
			3939: Pixel = 121;
			3940: Pixel = 121;
			3941: Pixel = 126;
			3942: Pixel = 112;
			3943: Pixel = 106;
			3944: Pixel = 109;
			3945: Pixel = 111;
			3946: Pixel = 113;
			3947: Pixel = 115;
			3948: Pixel = 120;
			3949: Pixel = 117;
			3950: Pixel = 117;
			3951: Pixel = 116;
			3952: Pixel = 113;
			3953: Pixel = 120;
			3954: Pixel = 125;
			3955: Pixel = 126;
			3956: Pixel = 128;
			3957: Pixel = 138;
			3958: Pixel = 135;
			3959: Pixel = 136;
			3960: Pixel = 137;
			3961: Pixel = 142;
			3962: Pixel = 142;
			3963: Pixel = 146;
			3964: Pixel = 146;
			3965: Pixel = 147;
			3966: Pixel = 156;
			3967: Pixel = 164;
			3968: Pixel = 175;
			3969: Pixel = 180;
			3970: Pixel = 180;
			3971: Pixel = 167;
			3972: Pixel = 162;
			3973: Pixel = 185;
			3974: Pixel = 206;
			3975: Pixel = 212;
			3976: Pixel = 207;
			3977: Pixel = 205;
			3978: Pixel = 204;
			3979: Pixel = 203;
			3980: Pixel = 208;
			3981: Pixel = 206;
			3982: Pixel = 203;
			3983: Pixel = 204;
			3984: Pixel = 207;
			3985: Pixel = 210;
			3986: Pixel = 213;
			3987: Pixel = 221;
			3988: Pixel = 232;
			3989: Pixel = 164;
			3990: Pixel = 72;
			3991: Pixel = 85;
			3992: Pixel = 91;
			3993: Pixel = 93;
			3994: Pixel = 94;
			3995: Pixel = 93;
			3996: Pixel = 97;
			3997: Pixel = 113;
			3998: Pixel = 131;
			3999: Pixel = 146;
			4000: Pixel = 155;
			4001: Pixel = 155;
			4002: Pixel = 154;
			4003: Pixel = 152;
			4004: Pixel = 151;
			4005: Pixel = 146;
			4006: Pixel = 130;
			4007: Pixel = 97;
			4008: Pixel = 51;
			4009: Pixel = 48;
			4010: Pixel = 87;
			4011: Pixel = 117;
			4012: Pixel = 136;
			4013: Pixel = 148;
			4014: Pixel = 148;
			4015: Pixel = 143;
			4016: Pixel = 145;
			4017: Pixel = 143;
			4018: Pixel = 142;
			4019: Pixel = 143;
			4020: Pixel = 144;
			4021: Pixel = 145;
			4022: Pixel = 144;
			4023: Pixel = 147;
			4024: Pixel = 151;
			4025: Pixel = 155;
			4026: Pixel = 91;
			4027: Pixel = 45;
			4028: Pixel = 58;
			4029: Pixel = 46;
			4030: Pixel = 46;
			4031: Pixel = 56;
			4032: Pixel = 53;
			4033: Pixel = 54;
			4034: Pixel = 53;
			4035: Pixel = 46;
			4036: Pixel = 47;
			4037: Pixel = 58;
			4038: Pixel = 51;
			4039: Pixel = 46;
			4040: Pixel = 48;
			4041: Pixel = 57;
			4042: Pixel = 66;
			4043: Pixel = 74;
			4044: Pixel = 79;
			4045: Pixel = 114;
			4046: Pixel = 146;
			4047: Pixel = 154;
			4048: Pixel = 140;
			4049: Pixel = 141;
			4050: Pixel = 119;
			4051: Pixel = 90;
			4052: Pixel = 84;
			4053: Pixel = 93;
			4054: Pixel = 90;
			4055: Pixel = 88;
			4056: Pixel = 85;
			4057: Pixel = 102;
			4058: Pixel = 131;
			4059: Pixel = 148;
			4060: Pixel = 159;
			4061: Pixel = 165;
			4062: Pixel = 168;
			4063: Pixel = 165;
			4064: Pixel = 164;
			4065: Pixel = 158;
			4066: Pixel = 146;
			4067: Pixel = 124;
			4068: Pixel = 99;
			4069: Pixel = 77;
			4070: Pixel = 81;
			4071: Pixel = 91;
			4072: Pixel = 97;
			4073: Pixel = 99;
			4074: Pixel = 97;
			4075: Pixel = 98;
			4076: Pixel = 99;
			4077: Pixel = 99;
			4078: Pixel = 99;
			4079: Pixel = 101;
			4080: Pixel = 104;
			4081: Pixel = 105;
			4082: Pixel = 111;
			4083: Pixel = 114;
			4084: Pixel = 116;
			4085: Pixel = 116;
			4086: Pixel = 118;
			4087: Pixel = 119;
			4088: Pixel = 121;
			4089: Pixel = 121;
			4090: Pixel = 125;
			4091: Pixel = 118;
			4092: Pixel = 106;
			4093: Pixel = 110;
			4094: Pixel = 114;
			4095: Pixel = 113;
			4096: Pixel = 114;
			4097: Pixel = 119;
			4098: Pixel = 118;
			4099: Pixel = 114;
			4100: Pixel = 112;
			4101: Pixel = 109;
			4102: Pixel = 116;
			4103: Pixel = 127;
			4104: Pixel = 129;
			4105: Pixel = 127;
			4106: Pixel = 134;
			4107: Pixel = 139;
			4108: Pixel = 139;
			4109: Pixel = 142;
			4110: Pixel = 143;
			4111: Pixel = 147;
			4112: Pixel = 140;
			4113: Pixel = 139;
			4114: Pixel = 141;
			4115: Pixel = 146;
			4116: Pixel = 156;
			4117: Pixel = 168;
			4118: Pixel = 179;
			4119: Pixel = 166;
			4120: Pixel = 151;
			4121: Pixel = 171;
			4122: Pixel = 204;
			4123: Pixel = 207;
			4124: Pixel = 201;
			4125: Pixel = 201;
			4126: Pixel = 206;
			4127: Pixel = 210;
			4128: Pixel = 205;
			4129: Pixel = 199;
			4130: Pixel = 197;
			4131: Pixel = 202;
			4132: Pixel = 203;
			4133: Pixel = 210;
			4134: Pixel = 212;
			4135: Pixel = 212;
			4136: Pixel = 212;
			4137: Pixel = 218;
			4138: Pixel = 223;
			4139: Pixel = 226;
			4140: Pixel = 126;
			4141: Pixel = 64;
			4142: Pixel = 79;
			4143: Pixel = 86;
			4144: Pixel = 88;
			4145: Pixel = 89;
			4146: Pixel = 96;
			4147: Pixel = 114;
			4148: Pixel = 133;
			4149: Pixel = 146;
			4150: Pixel = 155;
			4151: Pixel = 155;
			4152: Pixel = 153;
			4153: Pixel = 154;
			4154: Pixel = 153;
			4155: Pixel = 145;
			4156: Pixel = 131;
			4157: Pixel = 97;
			4158: Pixel = 49;
			4159: Pixel = 40;
			4160: Pixel = 73;
			4161: Pixel = 106;
			4162: Pixel = 127;
			4163: Pixel = 143;
			4164: Pixel = 149;
			4165: Pixel = 146;
			4166: Pixel = 144;
			4167: Pixel = 142;
			4168: Pixel = 142;
			4169: Pixel = 143;
			4170: Pixel = 143;
			4171: Pixel = 145;
			4172: Pixel = 145;
			4173: Pixel = 147;
			4174: Pixel = 159;
			4175: Pixel = 124;
			4176: Pixel = 44;
			4177: Pixel = 42;
			4178: Pixel = 48;
			4179: Pixel = 45;
			4180: Pixel = 51;
			4181: Pixel = 53;
			4182: Pixel = 52;
			4183: Pixel = 52;
			4184: Pixel = 45;
			4185: Pixel = 43;
			4186: Pixel = 57;
			4187: Pixel = 55;
			4188: Pixel = 46;
			4189: Pixel = 51;
			4190: Pixel = 50;
			4191: Pixel = 57;
			4192: Pixel = 70;
			4193: Pixel = 82;
			4194: Pixel = 112;
			4195: Pixel = 142;
			4196: Pixel = 148;
			4197: Pixel = 146;
			4198: Pixel = 140;
			4199: Pixel = 158;
			4200: Pixel = 96;
			4201: Pixel = 83;
			4202: Pixel = 87;
			4203: Pixel = 92;
			4204: Pixel = 91;
			4205: Pixel = 88;
			4206: Pixel = 85;
			4207: Pixel = 102;
			4208: Pixel = 130;
			4209: Pixel = 147;
			4210: Pixel = 158;
			4211: Pixel = 164;
			4212: Pixel = 167;
			4213: Pixel = 166;
			4214: Pixel = 163;
			4215: Pixel = 158;
			4216: Pixel = 145;
			4217: Pixel = 125;
			4218: Pixel = 101;
			4219: Pixel = 76;
			4220: Pixel = 79;
			4221: Pixel = 90;
			4222: Pixel = 96;
			4223: Pixel = 99;
			4224: Pixel = 99;
			4225: Pixel = 99;
			4226: Pixel = 99;
			4227: Pixel = 99;
			4228: Pixel = 101;
			4229: Pixel = 102;
			4230: Pixel = 104;
			4231: Pixel = 105;
			4232: Pixel = 110;
			4233: Pixel = 115;
			4234: Pixel = 119;
			4235: Pixel = 115;
			4236: Pixel = 117;
			4237: Pixel = 120;
			4238: Pixel = 120;
			4239: Pixel = 125;
			4240: Pixel = 125;
			4241: Pixel = 113;
			4242: Pixel = 113;
			4243: Pixel = 112;
			4244: Pixel = 112;
			4245: Pixel = 111;
			4246: Pixel = 116;
			4247: Pixel = 117;
			4248: Pixel = 114;
			4249: Pixel = 114;
			4250: Pixel = 114;
			4251: Pixel = 118;
			4252: Pixel = 121;
			4253: Pixel = 127;
			4254: Pixel = 129;
			4255: Pixel = 129;
			4256: Pixel = 136;
			4257: Pixel = 133;
			4258: Pixel = 136;
			4259: Pixel = 141;
			4260: Pixel = 145;
			4261: Pixel = 144;
			4262: Pixel = 137;
			4263: Pixel = 139;
			4264: Pixel = 142;
			4265: Pixel = 148;
			4266: Pixel = 159;
			4267: Pixel = 171;
			4268: Pixel = 147;
			4269: Pixel = 147;
			4270: Pixel = 182;
			4271: Pixel = 205;
			4272: Pixel = 202;
			4273: Pixel = 202;
			4274: Pixel = 203;
			4275: Pixel = 202;
			4276: Pixel = 203;
			4277: Pixel = 199;
			4278: Pixel = 195;
			4279: Pixel = 200;
			4280: Pixel = 201;
			4281: Pixel = 201;
			4282: Pixel = 202;
			4283: Pixel = 203;
			4284: Pixel = 202;
			4285: Pixel = 205;
			4286: Pixel = 207;
			4287: Pixel = 209;
			4288: Pixel = 212;
			4289: Pixel = 220;
			4290: Pixel = 212;
			4291: Pixel = 148;
			4292: Pixel = 81;
			4293: Pixel = 71;
			4294: Pixel = 83;
			4295: Pixel = 86;
			4296: Pixel = 92;
			4297: Pixel = 113;
			4298: Pixel = 133;
			4299: Pixel = 145;
			4300: Pixel = 154;
			4301: Pixel = 155;
			4302: Pixel = 154;
			4303: Pixel = 153;
			4304: Pixel = 152;
			4305: Pixel = 146;
			4306: Pixel = 131;
			4307: Pixel = 95;
			4308: Pixel = 50;
			4309: Pixel = 43;
			4310: Pixel = 58;
			4311: Pixel = 88;
			4312: Pixel = 117;
			4313: Pixel = 134;
			4314: Pixel = 146;
			4315: Pixel = 148;
			4316: Pixel = 144;
			4317: Pixel = 142;
			4318: Pixel = 141;
			4319: Pixel = 142;
			4320: Pixel = 144;
			4321: Pixel = 145;
			4322: Pixel = 147;
			4323: Pixel = 154;
			4324: Pixel = 146;
			4325: Pixel = 70;
			4326: Pixel = 36;
			4327: Pixel = 39;
			4328: Pixel = 43;
			4329: Pixel = 53;
			4330: Pixel = 57;
			4331: Pixel = 54;
			4332: Pixel = 53;
			4333: Pixel = 46;
			4334: Pixel = 41;
			4335: Pixel = 52;
			4336: Pixel = 57;
			4337: Pixel = 44;
			4338: Pixel = 51;
			4339: Pixel = 53;
			4340: Pixel = 57;
			4341: Pixel = 60;
			4342: Pixel = 68;
			4343: Pixel = 111;
			4344: Pixel = 140;
			4345: Pixel = 151;
			4346: Pixel = 145;
			4347: Pixel = 141;
			4348: Pixel = 157;
			4349: Pixel = 164;
			4350: Pixel = 86;
			4351: Pixel = 87;
			4352: Pixel = 90;
			4353: Pixel = 90;
			4354: Pixel = 91;
			4355: Pixel = 89;
			4356: Pixel = 85;
			4357: Pixel = 102;
			4358: Pixel = 128;
			4359: Pixel = 147;
			4360: Pixel = 158;
			4361: Pixel = 164;
			4362: Pixel = 165;
			4363: Pixel = 165;
			4364: Pixel = 164;
			4365: Pixel = 158;
			4366: Pixel = 144;
			4367: Pixel = 126;
			4368: Pixel = 101;
			4369: Pixel = 77;
			4370: Pixel = 76;
			4371: Pixel = 87;
			4372: Pixel = 94;
			4373: Pixel = 97;
			4374: Pixel = 100;
			4375: Pixel = 98;
			4376: Pixel = 99;
			4377: Pixel = 98;
			4378: Pixel = 101;
			4379: Pixel = 103;
			4380: Pixel = 103;
			4381: Pixel = 107;
			4382: Pixel = 110;
			4383: Pixel = 114;
			4384: Pixel = 116;
			4385: Pixel = 116;
			4386: Pixel = 117;
			4387: Pixel = 121;
			4388: Pixel = 118;
			4389: Pixel = 132;
			4390: Pixel = 118;
			4391: Pixel = 107;
			4392: Pixel = 112;
			4393: Pixel = 115;
			4394: Pixel = 110;
			4395: Pixel = 111;
			4396: Pixel = 114;
			4397: Pixel = 116;
			4398: Pixel = 115;
			4399: Pixel = 120;
			4400: Pixel = 120;
			4401: Pixel = 120;
			4402: Pixel = 129;
			4403: Pixel = 129;
			4404: Pixel = 128;
			4405: Pixel = 133;
			4406: Pixel = 140;
			4407: Pixel = 138;
			4408: Pixel = 137;
			4409: Pixel = 140;
			4410: Pixel = 139;
			4411: Pixel = 136;
			4412: Pixel = 133;
			4413: Pixel = 136;
			4414: Pixel = 142;
			4415: Pixel = 144;
			4416: Pixel = 155;
			4417: Pixel = 144;
			4418: Pixel = 156;
			4419: Pixel = 194;
			4420: Pixel = 195;
			4421: Pixel = 196;
			4422: Pixel = 199;
			4423: Pixel = 199;
			4424: Pixel = 205;
			4425: Pixel = 197;
			4426: Pixel = 199;
			4427: Pixel = 198;
			4428: Pixel = 195;
			4429: Pixel = 198;
			4430: Pixel = 201;
			4431: Pixel = 202;
			4432: Pixel = 202;
			4433: Pixel = 204;
			4434: Pixel = 204;
			4435: Pixel = 208;
			4436: Pixel = 210;
			4437: Pixel = 210;
			4438: Pixel = 210;
			4439: Pixel = 213;
			4440: Pixel = 219;
			4441: Pixel = 232;
			4442: Pixel = 181;
			4443: Pixel = 83;
			4444: Pixel = 69;
			4445: Pixel = 81;
			4446: Pixel = 89;
			4447: Pixel = 111;
			4448: Pixel = 132;
			4449: Pixel = 146;
			4450: Pixel = 154;
			4451: Pixel = 154;
			4452: Pixel = 154;
			4453: Pixel = 152;
			4454: Pixel = 156;
			4455: Pixel = 148;
			4456: Pixel = 128;
			4457: Pixel = 97;
			4458: Pixel = 55;
			4459: Pixel = 43;
			4460: Pixel = 41;
			4461: Pixel = 60;
			4462: Pixel = 97;
			4463: Pixel = 123;
			4464: Pixel = 139;
			4465: Pixel = 148;
			4466: Pixel = 146;
			4467: Pixel = 143;
			4468: Pixel = 140;
			4469: Pixel = 142;
			4470: Pixel = 144;
			4471: Pixel = 147;
			4472: Pixel = 151;
			4473: Pixel = 156;
			4474: Pixel = 96;
			4475: Pixel = 37;
			4476: Pixel = 39;
			4477: Pixel = 41;
			4478: Pixel = 47;
			4479: Pixel = 56;
			4480: Pixel = 56;
			4481: Pixel = 55;
			4482: Pixel = 52;
			4483: Pixel = 44;
			4484: Pixel = 48;
			4485: Pixel = 60;
			4486: Pixel = 49;
			4487: Pixel = 48;
			4488: Pixel = 52;
			4489: Pixel = 54;
			4490: Pixel = 55;
			4491: Pixel = 62;
			4492: Pixel = 95;
			4493: Pixel = 138;
			4494: Pixel = 145;
			4495: Pixel = 148;
			4496: Pixel = 143;
			4497: Pixel = 156;
			4498: Pixel = 166;
			4499: Pixel = 163;
			4500: Pixel = 86;
			4501: Pixel = 90;
			4502: Pixel = 93;
			4503: Pixel = 92;
			4504: Pixel = 93;
			4505: Pixel = 89;
			4506: Pixel = 89;
			4507: Pixel = 103;
			4508: Pixel = 130;
			4509: Pixel = 147;
			4510: Pixel = 158;
			4511: Pixel = 165;
			4512: Pixel = 166;
			4513: Pixel = 166;
			4514: Pixel = 163;
			4515: Pixel = 158;
			4516: Pixel = 146;
			4517: Pixel = 126;
			4518: Pixel = 102;
			4519: Pixel = 79;
			4520: Pixel = 76;
			4521: Pixel = 87;
			4522: Pixel = 93;
			4523: Pixel = 96;
			4524: Pixel = 96;
			4525: Pixel = 100;
			4526: Pixel = 101;
			4527: Pixel = 99;
			4528: Pixel = 100;
			4529: Pixel = 100;
			4530: Pixel = 102;
			4531: Pixel = 107;
			4532: Pixel = 109;
			4533: Pixel = 113;
			4534: Pixel = 117;
			4535: Pixel = 119;
			4536: Pixel = 119;
			4537: Pixel = 113;
			4538: Pixel = 131;
			4539: Pixel = 131;
			4540: Pixel = 105;
			4541: Pixel = 103;
			4542: Pixel = 105;
			4543: Pixel = 116;
			4544: Pixel = 115;
			4545: Pixel = 111;
			4546: Pixel = 113;
			4547: Pixel = 114;
			4548: Pixel = 113;
			4549: Pixel = 116;
			4550: Pixel = 118;
			4551: Pixel = 128;
			4552: Pixel = 132;
			4553: Pixel = 131;
			4554: Pixel = 137;
			4555: Pixel = 144;
			4556: Pixel = 139;
			4557: Pixel = 139;
			4558: Pixel = 141;
			4559: Pixel = 138;
			4560: Pixel = 137;
			4561: Pixel = 135;
			4562: Pixel = 133;
			4563: Pixel = 136;
			4564: Pixel = 139;
			4565: Pixel = 129;
			4566: Pixel = 139;
			4567: Pixel = 165;
			4568: Pixel = 196;
			4569: Pixel = 200;
			4570: Pixel = 195;
			4571: Pixel = 193;
			4572: Pixel = 192;
			4573: Pixel = 192;
			4574: Pixel = 193;
			4575: Pixel = 195;
			4576: Pixel = 195;
			4577: Pixel = 198;
			4578: Pixel = 200;
			4579: Pixel = 202;
			4580: Pixel = 203;
			4581: Pixel = 204;
			4582: Pixel = 208;
			4583: Pixel = 206;
			4584: Pixel = 207;
			4585: Pixel = 206;
			4586: Pixel = 205;
			4587: Pixel = 209;
			4588: Pixel = 207;
			4589: Pixel = 212;
			4590: Pixel = 211;
			4591: Pixel = 211;
			4592: Pixel = 232;
			4593: Pixel = 167;
			4594: Pixel = 57;
			4595: Pixel = 70;
			4596: Pixel = 86;
			4597: Pixel = 110;
			4598: Pixel = 131;
			4599: Pixel = 145;
			4600: Pixel = 154;
			4601: Pixel = 154;
			4602: Pixel = 153;
			4603: Pixel = 152;
			4604: Pixel = 154;
			4605: Pixel = 146;
			4606: Pixel = 128;
			4607: Pixel = 98;
			4608: Pixel = 57;
			4609: Pixel = 43;
			4610: Pixel = 40;
			4611: Pixel = 45;
			4612: Pixel = 72;
			4613: Pixel = 109;
			4614: Pixel = 132;
			4615: Pixel = 143;
			4616: Pixel = 148;
			4617: Pixel = 144;
			4618: Pixel = 140;
			4619: Pixel = 141;
			4620: Pixel = 146;
			4621: Pixel = 147;
			4622: Pixel = 156;
			4623: Pixel = 127;
			4624: Pixel = 48;
			4625: Pixel = 40;
			4626: Pixel = 44;
			4627: Pixel = 46;
			4628: Pixel = 51;
			4629: Pixel = 55;
			4630: Pixel = 52;
			4631: Pixel = 56;
			4632: Pixel = 49;
			4633: Pixel = 46;
			4634: Pixel = 55;
			4635: Pixel = 49;
			4636: Pixel = 44;
			4637: Pixel = 53;
			4638: Pixel = 55;
			4639: Pixel = 51;
			4640: Pixel = 51;
			4641: Pixel = 87;
			4642: Pixel = 138;
			4643: Pixel = 145;
			4644: Pixel = 141;
			4645: Pixel = 139;
			4646: Pixel = 150;
			4647: Pixel = 165;
			4648: Pixel = 164;
			4649: Pixel = 162;
			4650: Pixel = 87;
			4651: Pixel = 90;
			4652: Pixel = 93;
			4653: Pixel = 91;
			4654: Pixel = 91;
			4655: Pixel = 90;
			4656: Pixel = 89;
			4657: Pixel = 105;
			4658: Pixel = 130;
			4659: Pixel = 147;
			4660: Pixel = 158;
			4661: Pixel = 163;
			4662: Pixel = 163;
			4663: Pixel = 163;
			4664: Pixel = 162;
			4665: Pixel = 159;
			4666: Pixel = 147;
			4667: Pixel = 127;
			4668: Pixel = 100;
			4669: Pixel = 79;
			4670: Pixel = 77;
			4671: Pixel = 87;
			4672: Pixel = 93;
			4673: Pixel = 95;
			4674: Pixel = 97;
			4675: Pixel = 100;
			4676: Pixel = 101;
			4677: Pixel = 99;
			4678: Pixel = 97;
			4679: Pixel = 100;
			4680: Pixel = 102;
			4681: Pixel = 106;
			4682: Pixel = 110;
			4683: Pixel = 114;
			4684: Pixel = 115;
			4685: Pixel = 116;
			4686: Pixel = 115;
			4687: Pixel = 109;
			4688: Pixel = 165;
			4689: Pixel = 124;
			4690: Pixel = 97;
			4691: Pixel = 106;
			4692: Pixel = 107;
			4693: Pixel = 112;
			4694: Pixel = 113;
			4695: Pixel = 112;
			4696: Pixel = 113;
			4697: Pixel = 113;
			4698: Pixel = 113;
			4699: Pixel = 119;
			4700: Pixel = 124;
			4701: Pixel = 122;
			4702: Pixel = 131;
			4703: Pixel = 134;
			4704: Pixel = 144;
			4705: Pixel = 139;
			4706: Pixel = 130;
			4707: Pixel = 137;
			4708: Pixel = 142;
			4709: Pixel = 140;
			4710: Pixel = 136;
			4711: Pixel = 131;
			4712: Pixel = 128;
			4713: Pixel = 126;
			4714: Pixel = 123;
			4715: Pixel = 149;
			4716: Pixel = 186;
			4717: Pixel = 183;
			4718: Pixel = 189;
			4719: Pixel = 197;
			4720: Pixel = 192;
			4721: Pixel = 191;
			4722: Pixel = 191;
			4723: Pixel = 189;
			4724: Pixel = 187;
			4725: Pixel = 187;
			4726: Pixel = 195;
			4727: Pixel = 202;
			4728: Pixel = 206;
			4729: Pixel = 202;
			4730: Pixel = 205;
			4731: Pixel = 204;
			4732: Pixel = 202;
			4733: Pixel = 206;
			4734: Pixel = 206;
			4735: Pixel = 208;
			4736: Pixel = 206;
			4737: Pixel = 206;
			4738: Pixel = 204;
			4739: Pixel = 206;
			4740: Pixel = 213;
			4741: Pixel = 215;
			4742: Pixel = 217;
			4743: Pixel = 226;
			4744: Pixel = 111;
			4745: Pixel = 59;
			4746: Pixel = 81;
			4747: Pixel = 105;
			4748: Pixel = 128;
			4749: Pixel = 144;
			4750: Pixel = 152;
			4751: Pixel = 154;
			4752: Pixel = 155;
			4753: Pixel = 153;
			4754: Pixel = 152;
			4755: Pixel = 146;
			4756: Pixel = 130;
			4757: Pixel = 101;
			4758: Pixel = 58;
			4759: Pixel = 43;
			4760: Pixel = 45;
			4761: Pixel = 39;
			4762: Pixel = 48;
			4763: Pixel = 84;
			4764: Pixel = 118;
			4765: Pixel = 132;
			4766: Pixel = 139;
			4767: Pixel = 138;
			4768: Pixel = 134;
			4769: Pixel = 138;
			4770: Pixel = 142;
			4771: Pixel = 152;
			4772: Pixel = 148;
			4773: Pixel = 71;
			4774: Pixel = 39;
			4775: Pixel = 44;
			4776: Pixel = 46;
			4777: Pixel = 49;
			4778: Pixel = 53;
			4779: Pixel = 54;
			4780: Pixel = 55;
			4781: Pixel = 52;
			4782: Pixel = 46;
			4783: Pixel = 52;
			4784: Pixel = 55;
			4785: Pixel = 45;
			4786: Pixel = 52;
			4787: Pixel = 54;
			4788: Pixel = 49;
			4789: Pixel = 46;
			4790: Pixel = 74;
			4791: Pixel = 129;
			4792: Pixel = 153;
			4793: Pixel = 142;
			4794: Pixel = 133;
			4795: Pixel = 147;
			4796: Pixel = 161;
			4797: Pixel = 163;
			4798: Pixel = 163;
			4799: Pixel = 164;
			4800: Pixel = 92;
			4801: Pixel = 91;
			4802: Pixel = 92;
			4803: Pixel = 91;
			4804: Pixel = 92;
			4805: Pixel = 89;
			4806: Pixel = 85;
			4807: Pixel = 101;
			4808: Pixel = 130;
			4809: Pixel = 148;
			4810: Pixel = 158;
			4811: Pixel = 163;
			4812: Pixel = 165;
			4813: Pixel = 163;
			4814: Pixel = 163;
			4815: Pixel = 162;
			4816: Pixel = 148;
			4817: Pixel = 127;
			4818: Pixel = 101;
			4819: Pixel = 77;
			4820: Pixel = 79;
			4821: Pixel = 86;
			4822: Pixel = 91;
			4823: Pixel = 96;
			4824: Pixel = 97;
			4825: Pixel = 98;
			4826: Pixel = 101;
			4827: Pixel = 102;
			4828: Pixel = 100;
			4829: Pixel = 102;
			4830: Pixel = 106;
			4831: Pixel = 108;
			4832: Pixel = 111;
			4833: Pixel = 113;
			4834: Pixel = 114;
			4835: Pixel = 115;
			4836: Pixel = 106;
			4837: Pixel = 126;
			4838: Pixel = 182;
			4839: Pixel = 107;
			4840: Pixel = 101;
			4841: Pixel = 107;
			4842: Pixel = 108;
			4843: Pixel = 109;
			4844: Pixel = 110;
			4845: Pixel = 113;
			4846: Pixel = 115;
			4847: Pixel = 119;
			4848: Pixel = 120;
			4849: Pixel = 121;
			4850: Pixel = 126;
			4851: Pixel = 125;
			4852: Pixel = 133;
			4853: Pixel = 140;
			4854: Pixel = 136;
			4855: Pixel = 130;
			4856: Pixel = 133;
			4857: Pixel = 136;
			4858: Pixel = 140;
			4859: Pixel = 137;
			4860: Pixel = 129;
			4861: Pixel = 128;
			4862: Pixel = 110;
			4863: Pixel = 123;
			4864: Pixel = 160;
			4865: Pixel = 180;
			4866: Pixel = 192;
			4867: Pixel = 193;
			4868: Pixel = 183;
			4869: Pixel = 185;
			4870: Pixel = 192;
			4871: Pixel = 190;
			4872: Pixel = 181;
			4873: Pixel = 190;
			4874: Pixel = 194;
			4875: Pixel = 196;
			4876: Pixel = 197;
			4877: Pixel = 199;
			4878: Pixel = 202;
			4879: Pixel = 206;
			4880: Pixel = 202;
			4881: Pixel = 204;
			4882: Pixel = 203;
			4883: Pixel = 206;
			4884: Pixel = 203;
			4885: Pixel = 200;
			4886: Pixel = 202;
			4887: Pixel = 205;
			4888: Pixel = 205;
			4889: Pixel = 204;
			4890: Pixel = 212;
			4891: Pixel = 214;
			4892: Pixel = 217;
			4893: Pixel = 228;
			4894: Pixel = 203;
			4895: Pixel = 83;
			4896: Pixel = 67;
			4897: Pixel = 102;
			4898: Pixel = 129;
			4899: Pixel = 143;
			4900: Pixel = 151;
			4901: Pixel = 152;
			4902: Pixel = 154;
			4903: Pixel = 153;
			4904: Pixel = 154;
			4905: Pixel = 145;
			4906: Pixel = 128;
			4907: Pixel = 100;
			4908: Pixel = 62;
			4909: Pixel = 45;
			4910: Pixel = 45;
			4911: Pixel = 42;
			4912: Pixel = 40;
			4913: Pixel = 53;
			4914: Pixel = 80;
			4915: Pixel = 114;
			4916: Pixel = 157;
			4917: Pixel = 180;
			4918: Pixel = 165;
			4919: Pixel = 143;
			4920: Pixel = 157;
			4921: Pixel = 149;
			4922: Pixel = 99;
			4923: Pixel = 40;
			4924: Pixel = 44;
			4925: Pixel = 46;
			4926: Pixel = 49;
			4927: Pixel = 55;
			4928: Pixel = 53;
			4929: Pixel = 52;
			4930: Pixel = 55;
			4931: Pixel = 51;
			4932: Pixel = 50;
			4933: Pixel = 55;
			4934: Pixel = 48;
			4935: Pixel = 50;
			4936: Pixel = 56;
			4937: Pixel = 52;
			4938: Pixel = 37;
			4939: Pixel = 54;
			4940: Pixel = 119;
			4941: Pixel = 152;
			4942: Pixel = 145;
			4943: Pixel = 134;
			4944: Pixel = 144;
			4945: Pixel = 159;
			4946: Pixel = 161;
			4947: Pixel = 161;
			4948: Pixel = 160;
			4949: Pixel = 161;
			4950: Pixel = 92;
			4951: Pixel = 91;
			4952: Pixel = 90;
			4953: Pixel = 89;
			4954: Pixel = 89;
			4955: Pixel = 87;
			4956: Pixel = 84;
			4957: Pixel = 99;
			4958: Pixel = 129;
			4959: Pixel = 147;
			4960: Pixel = 157;
			4961: Pixel = 164;
			4962: Pixel = 164;
			4963: Pixel = 163;
			4964: Pixel = 163;
			4965: Pixel = 161;
			4966: Pixel = 147;
			4967: Pixel = 129;
			4968: Pixel = 104;
			4969: Pixel = 78;
			4970: Pixel = 77;
			4971: Pixel = 86;
			4972: Pixel = 93;
			4973: Pixel = 93;
			4974: Pixel = 94;
			4975: Pixel = 98;
			4976: Pixel = 100;
			4977: Pixel = 100;
			4978: Pixel = 99;
			4979: Pixel = 104;
			4980: Pixel = 107;
			4981: Pixel = 107;
			4982: Pixel = 109;
			4983: Pixel = 112;
			4984: Pixel = 114;
			4985: Pixel = 112;
			4986: Pixel = 98;
			4987: Pixel = 165;
			4988: Pixel = 175;
			4989: Pixel = 97;
			4990: Pixel = 105;
			4991: Pixel = 103;
			4992: Pixel = 107;
			4993: Pixel = 111;
			4994: Pixel = 113;
			4995: Pixel = 111;
			4996: Pixel = 109;
			4997: Pixel = 117;
			4998: Pixel = 119;
			4999: Pixel = 123;
			5000: Pixel = 128;
			5001: Pixel = 132;
			5002: Pixel = 134;
			5003: Pixel = 135;
			5004: Pixel = 138;
			5005: Pixel = 134;
			5006: Pixel = 132;
			5007: Pixel = 139;
			5008: Pixel = 137;
			5009: Pixel = 125;
			5010: Pixel = 123;
			5011: Pixel = 111;
			5012: Pixel = 129;
			5013: Pixel = 167;
			5014: Pixel = 190;
			5015: Pixel = 187;
			5016: Pixel = 183;
			5017: Pixel = 184;
			5018: Pixel = 190;
			5019: Pixel = 187;
			5020: Pixel = 175;
			5021: Pixel = 177;
			5022: Pixel = 187;
			5023: Pixel = 196;
			5024: Pixel = 198;
			5025: Pixel = 197;
			5026: Pixel = 195;
			5027: Pixel = 196;
			5028: Pixel = 201;
			5029: Pixel = 204;
			5030: Pixel = 202;
			5031: Pixel = 201;
			5032: Pixel = 202;
			5033: Pixel = 200;
			5034: Pixel = 201;
			5035: Pixel = 199;
			5036: Pixel = 201;
			5037: Pixel = 207;
			5038: Pixel = 210;
			5039: Pixel = 205;
			5040: Pixel = 207;
			5041: Pixel = 211;
			5042: Pixel = 213;
			5043: Pixel = 220;
			5044: Pixel = 238;
			5045: Pixel = 144;
			5046: Pixel = 53;
			5047: Pixel = 101;
			5048: Pixel = 128;
			5049: Pixel = 144;
			5050: Pixel = 151;
			5051: Pixel = 151;
			5052: Pixel = 153;
			5053: Pixel = 153;
			5054: Pixel = 154;
			5055: Pixel = 148;
			5056: Pixel = 130;
			5057: Pixel = 101;
			5058: Pixel = 61;
			5059: Pixel = 44;
			5060: Pixel = 45;
			5061: Pixel = 45;
			5062: Pixel = 39;
			5063: Pixel = 27;
			5064: Pixel = 95;
			5065: Pixel = 194;
			5066: Pixel = 217;
			5067: Pixel = 210;
			5068: Pixel = 203;
			5069: Pixel = 201;
			5070: Pixel = 216;
			5071: Pixel = 153;
			5072: Pixel = 45;
			5073: Pixel = 42;
			5074: Pixel = 47;
			5075: Pixel = 47;
			5076: Pixel = 53;
			5077: Pixel = 55;
			5078: Pixel = 53;
			5079: Pixel = 54;
			5080: Pixel = 58;
			5081: Pixel = 53;
			5082: Pixel = 54;
			5083: Pixel = 48;
			5084: Pixel = 48;
			5085: Pixel = 57;
			5086: Pixel = 50;
			5087: Pixel = 43;
			5088: Pixel = 51;
			5089: Pixel = 101;
			5090: Pixel = 148;
			5091: Pixel = 148;
			5092: Pixel = 136;
			5093: Pixel = 141;
			5094: Pixel = 158;
			5095: Pixel = 162;
			5096: Pixel = 160;
			5097: Pixel = 159;
			5098: Pixel = 158;
			5099: Pixel = 158;
			5100: Pixel = 89;
			5101: Pixel = 89;
			5102: Pixel = 89;
			5103: Pixel = 87;
			5104: Pixel = 90;
			5105: Pixel = 88;
			5106: Pixel = 82;
			5107: Pixel = 97;
			5108: Pixel = 127;
			5109: Pixel = 146;
			5110: Pixel = 159;
			5111: Pixel = 164;
			5112: Pixel = 163;
			5113: Pixel = 163;
			5114: Pixel = 163;
			5115: Pixel = 159;
			5116: Pixel = 146;
			5117: Pixel = 127;
			5118: Pixel = 100;
			5119: Pixel = 73;
			5120: Pixel = 75;
			5121: Pixel = 84;
			5122: Pixel = 88;
			5123: Pixel = 91;
			5124: Pixel = 95;
			5125: Pixel = 95;
			5126: Pixel = 96;
			5127: Pixel = 95;
			5128: Pixel = 98;
			5129: Pixel = 100;
			5130: Pixel = 102;
			5131: Pixel = 105;
			5132: Pixel = 107;
			5133: Pixel = 109;
			5134: Pixel = 111;
			5135: Pixel = 105;
			5136: Pixel = 105;
			5137: Pixel = 197;
			5138: Pixel = 152;
			5139: Pixel = 98;
			5140: Pixel = 102;
			5141: Pixel = 105;
			5142: Pixel = 108;
			5143: Pixel = 113;
			5144: Pixel = 113;
			5145: Pixel = 113;
			5146: Pixel = 113;
			5147: Pixel = 118;
			5148: Pixel = 118;
			5149: Pixel = 125;
			5150: Pixel = 130;
			5151: Pixel = 135;
			5152: Pixel = 137;
			5153: Pixel = 133;
			5154: Pixel = 132;
			5155: Pixel = 129;
			5156: Pixel = 137;
			5157: Pixel = 133;
			5158: Pixel = 119;
			5159: Pixel = 107;
			5160: Pixel = 115;
			5161: Pixel = 143;
			5162: Pixel = 175;
			5163: Pixel = 178;
			5164: Pixel = 190;
			5165: Pixel = 182;
			5166: Pixel = 173;
			5167: Pixel = 176;
			5168: Pixel = 184;
			5169: Pixel = 181;
			5170: Pixel = 183;
			5171: Pixel = 187;
			5172: Pixel = 188;
			5173: Pixel = 193;
			5174: Pixel = 196;
			5175: Pixel = 195;
			5176: Pixel = 195;
			5177: Pixel = 196;
			5178: Pixel = 196;
			5179: Pixel = 199;
			5180: Pixel = 198;
			5181: Pixel = 193;
			5182: Pixel = 196;
			5183: Pixel = 203;
			5184: Pixel = 204;
			5185: Pixel = 207;
			5186: Pixel = 202;
			5187: Pixel = 204;
			5188: Pixel = 207;
			5189: Pixel = 207;
			5190: Pixel = 207;
			5191: Pixel = 208;
			5192: Pixel = 210;
			5193: Pixel = 215;
			5194: Pixel = 229;
			5195: Pixel = 195;
			5196: Pixel = 67;
			5197: Pixel = 89;
			5198: Pixel = 126;
			5199: Pixel = 143;
			5200: Pixel = 150;
			5201: Pixel = 153;
			5202: Pixel = 153;
			5203: Pixel = 154;
			5204: Pixel = 153;
			5205: Pixel = 148;
			5206: Pixel = 128;
			5207: Pixel = 100;
			5208: Pixel = 60;
			5209: Pixel = 43;
			5210: Pixel = 45;
			5211: Pixel = 35;
			5212: Pixel = 32;
			5213: Pixel = 110;
			5214: Pixel = 215;
			5215: Pixel = 211;
			5216: Pixel = 194;
			5217: Pixel = 201;
			5218: Pixel = 216;
			5219: Pixel = 224;
			5220: Pixel = 229;
			5221: Pixel = 202;
			5222: Pixel = 53;
			5223: Pixel = 40;
			5224: Pixel = 46;
			5225: Pixel = 48;
			5226: Pixel = 57;
			5227: Pixel = 52;
			5228: Pixel = 58;
			5229: Pixel = 54;
			5230: Pixel = 50;
			5231: Pixel = 52;
			5232: Pixel = 54;
			5233: Pixel = 49;
			5234: Pixel = 53;
			5235: Pixel = 59;
			5236: Pixel = 47;
			5237: Pixel = 38;
			5238: Pixel = 84;
			5239: Pixel = 143;
			5240: Pixel = 151;
			5241: Pixel = 141;
			5242: Pixel = 141;
			5243: Pixel = 157;
			5244: Pixel = 164;
			5245: Pixel = 161;
			5246: Pixel = 159;
			5247: Pixel = 159;
			5248: Pixel = 157;
			5249: Pixel = 158;
			5250: Pixel = 88;
			5251: Pixel = 89;
			5252: Pixel = 90;
			5253: Pixel = 91;
			5254: Pixel = 93;
			5255: Pixel = 91;
			5256: Pixel = 85;
			5257: Pixel = 99;
			5258: Pixel = 127;
			5259: Pixel = 144;
			5260: Pixel = 158;
			5261: Pixel = 163;
			5262: Pixel = 165;
			5263: Pixel = 164;
			5264: Pixel = 163;
			5265: Pixel = 160;
			5266: Pixel = 146;
			5267: Pixel = 127;
			5268: Pixel = 97;
			5269: Pixel = 71;
			5270: Pixel = 73;
			5271: Pixel = 80;
			5272: Pixel = 89;
			5273: Pixel = 93;
			5274: Pixel = 97;
			5275: Pixel = 98;
			5276: Pixel = 98;
			5277: Pixel = 97;
			5278: Pixel = 98;
			5279: Pixel = 99;
			5280: Pixel = 104;
			5281: Pixel = 105;
			5282: Pixel = 105;
			5283: Pixel = 111;
			5284: Pixel = 112;
			5285: Pixel = 99;
			5286: Pixel = 131;
			5287: Pixel = 206;
			5288: Pixel = 146;
			5289: Pixel = 102;
			5290: Pixel = 100;
			5291: Pixel = 106;
			5292: Pixel = 108;
			5293: Pixel = 109;
			5294: Pixel = 116;
			5295: Pixel = 114;
			5296: Pixel = 118;
			5297: Pixel = 116;
			5298: Pixel = 121;
			5299: Pixel = 129;
			5300: Pixel = 129;
			5301: Pixel = 126;
			5302: Pixel = 126;
			5303: Pixel = 118;
			5304: Pixel = 131;
			5305: Pixel = 137;
			5306: Pixel = 131;
			5307: Pixel = 125;
			5308: Pixel = 111;
			5309: Pixel = 114;
			5310: Pixel = 156;
			5311: Pixel = 178;
			5312: Pixel = 181;
			5313: Pixel = 174;
			5314: Pixel = 167;
			5315: Pixel = 177;
			5316: Pixel = 180;
			5317: Pixel = 172;
			5318: Pixel = 169;
			5319: Pixel = 182;
			5320: Pixel = 187;
			5321: Pixel = 186;
			5322: Pixel = 186;
			5323: Pixel = 193;
			5324: Pixel = 192;
			5325: Pixel = 195;
			5326: Pixel = 195;
			5327: Pixel = 193;
			5328: Pixel = 189;
			5329: Pixel = 189;
			5330: Pixel = 193;
			5331: Pixel = 201;
			5332: Pixel = 203;
			5333: Pixel = 203;
			5334: Pixel = 204;
			5335: Pixel = 199;
			5336: Pixel = 203;
			5337: Pixel = 199;
			5338: Pixel = 203;
			5339: Pixel = 205;
			5340: Pixel = 205;
			5341: Pixel = 203;
			5342: Pixel = 205;
			5343: Pixel = 208;
			5344: Pixel = 219;
			5345: Pixel = 229;
			5346: Pixel = 129;
			5347: Pixel = 74;
			5348: Pixel = 124;
			5349: Pixel = 143;
			5350: Pixel = 152;
			5351: Pixel = 153;
			5352: Pixel = 155;
			5353: Pixel = 154;
			5354: Pixel = 153;
			5355: Pixel = 148;
			5356: Pixel = 128;
			5357: Pixel = 96;
			5358: Pixel = 55;
			5359: Pixel = 41;
			5360: Pixel = 32;
			5361: Pixel = 43;
			5362: Pixel = 145;
			5363: Pixel = 221;
			5364: Pixel = 192;
			5365: Pixel = 184;
			5366: Pixel = 213;
			5367: Pixel = 221;
			5368: Pixel = 223;
			5369: Pixel = 223;
			5370: Pixel = 227;
			5371: Pixel = 239;
			5372: Pixel = 104;
			5373: Pixel = 32;
			5374: Pixel = 46;
			5375: Pixel = 48;
			5376: Pixel = 54;
			5377: Pixel = 55;
			5378: Pixel = 52;
			5379: Pixel = 49;
			5380: Pixel = 49;
			5381: Pixel = 52;
			5382: Pixel = 47;
			5383: Pixel = 50;
			5384: Pixel = 54;
			5385: Pixel = 53;
			5386: Pixel = 45;
			5387: Pixel = 65;
			5388: Pixel = 128;
			5389: Pixel = 153;
			5390: Pixel = 144;
			5391: Pixel = 140;
			5392: Pixel = 153;
			5393: Pixel = 161;
			5394: Pixel = 161;
			5395: Pixel = 160;
			5396: Pixel = 159;
			5397: Pixel = 158;
			5398: Pixel = 158;
			5399: Pixel = 157;
			5400: Pixel = 91;
			5401: Pixel = 91;
			5402: Pixel = 92;
			5403: Pixel = 93;
			5404: Pixel = 96;
			5405: Pixel = 93;
			5406: Pixel = 86;
			5407: Pixel = 99;
			5408: Pixel = 125;
			5409: Pixel = 145;
			5410: Pixel = 157;
			5411: Pixel = 166;
			5412: Pixel = 167;
			5413: Pixel = 166;
			5414: Pixel = 164;
			5415: Pixel = 159;
			5416: Pixel = 146;
			5417: Pixel = 126;
			5418: Pixel = 96;
			5419: Pixel = 74;
			5420: Pixel = 74;
			5421: Pixel = 78;
			5422: Pixel = 90;
			5423: Pixel = 95;
			5424: Pixel = 99;
			5425: Pixel = 98;
			5426: Pixel = 100;
			5427: Pixel = 100;
			5428: Pixel = 100;
			5429: Pixel = 99;
			5430: Pixel = 102;
			5431: Pixel = 105;
			5432: Pixel = 108;
			5433: Pixel = 112;
			5434: Pixel = 116;
			5435: Pixel = 99;
			5436: Pixel = 160;
			5437: Pixel = 205;
			5438: Pixel = 131;
			5439: Pixel = 96;
			5440: Pixel = 101;
			5441: Pixel = 104;
			5442: Pixel = 106;
			5443: Pixel = 116;
			5444: Pixel = 110;
			5445: Pixel = 111;
			5446: Pixel = 115;
			5447: Pixel = 119;
			5448: Pixel = 129;
			5449: Pixel = 130;
			5450: Pixel = 122;
			5451: Pixel = 118;
			5452: Pixel = 119;
			5453: Pixel = 130;
			5454: Pixel = 131;
			5455: Pixel = 128;
			5456: Pixel = 121;
			5457: Pixel = 105;
			5458: Pixel = 119;
			5459: Pixel = 166;
			5460: Pixel = 175;
			5461: Pixel = 179;
			5462: Pixel = 169;
			5463: Pixel = 164;
			5464: Pixel = 166;
			5465: Pixel = 173;
			5466: Pixel = 171;
			5467: Pixel = 181;
			5468: Pixel = 183;
			5469: Pixel = 171;
			5470: Pixel = 184;
			5471: Pixel = 193;
			5472: Pixel = 188;
			5473: Pixel = 187;
			5474: Pixel = 188;
			5475: Pixel = 192;
			5476: Pixel = 193;
			5477: Pixel = 184;
			5478: Pixel = 189;
			5479: Pixel = 194;
			5480: Pixel = 200;
			5481: Pixel = 199;
			5482: Pixel = 195;
			5483: Pixel = 202;
			5484: Pixel = 200;
			5485: Pixel = 200;
			5486: Pixel = 198;
			5487: Pixel = 198;
			5488: Pixel = 202;
			5489: Pixel = 207;
			5490: Pixel = 205;
			5491: Pixel = 207;
			5492: Pixel = 207;
			5493: Pixel = 206;
			5494: Pixel = 210;
			5495: Pixel = 223;
			5496: Pixel = 206;
			5497: Pixel = 93;
			5498: Pixel = 112;
			5499: Pixel = 141;
			5500: Pixel = 155;
			5501: Pixel = 155;
			5502: Pixel = 157;
			5503: Pixel = 155;
			5504: Pixel = 154;
			5505: Pixel = 146;
			5506: Pixel = 126;
			5507: Pixel = 91;
			5508: Pixel = 44;
			5509: Pixel = 24;
			5510: Pixel = 63;
			5511: Pixel = 178;
			5512: Pixel = 218;
			5513: Pixel = 174;
			5514: Pixel = 184;
			5515: Pixel = 220;
			5516: Pixel = 217;
			5517: Pixel = 213;
			5518: Pixel = 214;
			5519: Pixel = 210;
			5520: Pixel = 214;
			5521: Pixel = 240;
			5522: Pixel = 143;
			5523: Pixel = 31;
			5524: Pixel = 46;
			5525: Pixel = 49;
			5526: Pixel = 51;
			5527: Pixel = 55;
			5528: Pixel = 51;
			5529: Pixel = 48;
			5530: Pixel = 50;
			5531: Pixel = 44;
			5532: Pixel = 47;
			5533: Pixel = 52;
			5534: Pixel = 56;
			5535: Pixel = 51;
			5536: Pixel = 51;
			5537: Pixel = 108;
			5538: Pixel = 153;
			5539: Pixel = 148;
			5540: Pixel = 140;
			5541: Pixel = 150;
			5542: Pixel = 160;
			5543: Pixel = 159;
			5544: Pixel = 158;
			5545: Pixel = 159;
			5546: Pixel = 158;
			5547: Pixel = 158;
			5548: Pixel = 157;
			5549: Pixel = 157;
			5550: Pixel = 92;
			5551: Pixel = 93;
			5552: Pixel = 94;
			5553: Pixel = 96;
			5554: Pixel = 96;
			5555: Pixel = 97;
			5556: Pixel = 93;
			5557: Pixel = 101;
			5558: Pixel = 126;
			5559: Pixel = 144;
			5560: Pixel = 158;
			5561: Pixel = 167;
			5562: Pixel = 167;
			5563: Pixel = 167;
			5564: Pixel = 166;
			5565: Pixel = 159;
			5566: Pixel = 148;
			5567: Pixel = 127;
			5568: Pixel = 98;
			5569: Pixel = 75;
			5570: Pixel = 76;
			5571: Pixel = 82;
			5572: Pixel = 91;
			5573: Pixel = 96;
			5574: Pixel = 99;
			5575: Pixel = 98;
			5576: Pixel = 101;
			5577: Pixel = 100;
			5578: Pixel = 100;
			5579: Pixel = 103;
			5580: Pixel = 104;
			5581: Pixel = 106;
			5582: Pixel = 110;
			5583: Pixel = 112;
			5584: Pixel = 112;
			5585: Pixel = 99;
			5586: Pixel = 181;
			5587: Pixel = 196;
			5588: Pixel = 132;
			5589: Pixel = 93;
			5590: Pixel = 102;
			5591: Pixel = 105;
			5592: Pixel = 109;
			5593: Pixel = 103;
			5594: Pixel = 102;
			5595: Pixel = 116;
			5596: Pixel = 120;
			5597: Pixel = 127;
			5598: Pixel = 125;
			5599: Pixel = 121;
			5600: Pixel = 115;
			5601: Pixel = 122;
			5602: Pixel = 137;
			5603: Pixel = 128;
			5604: Pixel = 127;
			5605: Pixel = 127;
			5606: Pixel = 104;
			5607: Pixel = 127;
			5608: Pixel = 160;
			5609: Pixel = 174;
			5610: Pixel = 176;
			5611: Pixel = 162;
			5612: Pixel = 160;
			5613: Pixel = 173;
			5614: Pixel = 170;
			5615: Pixel = 175;
			5616: Pixel = 181;
			5617: Pixel = 175;
			5618: Pixel = 179;
			5619: Pixel = 185;
			5620: Pixel = 186;
			5621: Pixel = 187;
			5622: Pixel = 188;
			5623: Pixel = 186;
			5624: Pixel = 185;
			5625: Pixel = 180;
			5626: Pixel = 179;
			5627: Pixel = 189;
			5628: Pixel = 200;
			5629: Pixel = 200;
			5630: Pixel = 194;
			5631: Pixel = 196;
			5632: Pixel = 193;
			5633: Pixel = 193;
			5634: Pixel = 202;
			5635: Pixel = 199;
			5636: Pixel = 201;
			5637: Pixel = 207;
			5638: Pixel = 202;
			5639: Pixel = 201;
			5640: Pixel = 199;
			5641: Pixel = 203;
			5642: Pixel = 203;
			5643: Pixel = 205;
			5644: Pixel = 206;
			5645: Pixel = 208;
			5646: Pixel = 222;
			5647: Pixel = 165;
			5648: Pixel = 107;
			5649: Pixel = 138;
			5650: Pixel = 152;
			5651: Pixel = 155;
			5652: Pixel = 156;
			5653: Pixel = 155;
			5654: Pixel = 152;
			5655: Pixel = 142;
			5656: Pixel = 118;
			5657: Pixel = 73;
			5658: Pixel = 35;
			5659: Pixel = 97;
			5660: Pixel = 202;
			5661: Pixel = 211;
			5662: Pixel = 168;
			5663: Pixel = 192;
			5664: Pixel = 219;
			5665: Pixel = 215;
			5666: Pixel = 209;
			5667: Pixel = 203;
			5668: Pixel = 206;
			5669: Pixel = 205;
			5670: Pixel = 213;
			5671: Pixel = 238;
			5672: Pixel = 155;
			5673: Pixel = 30;
			5674: Pixel = 46;
			5675: Pixel = 51;
			5676: Pixel = 53;
			5677: Pixel = 50;
			5678: Pixel = 45;
			5679: Pixel = 47;
			5680: Pixel = 46;
			5681: Pixel = 43;
			5682: Pixel = 49;
			5683: Pixel = 53;
			5684: Pixel = 51;
			5685: Pixel = 42;
			5686: Pixel = 79;
			5687: Pixel = 146;
			5688: Pixel = 155;
			5689: Pixel = 143;
			5690: Pixel = 147;
			5691: Pixel = 159;
			5692: Pixel = 160;
			5693: Pixel = 157;
			5694: Pixel = 157;
			5695: Pixel = 158;
			5696: Pixel = 157;
			5697: Pixel = 156;
			5698: Pixel = 157;
			5699: Pixel = 158;
			5700: Pixel = 95;
			5701: Pixel = 96;
			5702: Pixel = 97;
			5703: Pixel = 100;
			5704: Pixel = 98;
			5705: Pixel = 97;
			5706: Pixel = 94;
			5707: Pixel = 101;
			5708: Pixel = 126;
			5709: Pixel = 145;
			5710: Pixel = 158;
			5711: Pixel = 166;
			5712: Pixel = 167;
			5713: Pixel = 167;
			5714: Pixel = 166;
			5715: Pixel = 163;
			5716: Pixel = 152;
			5717: Pixel = 129;
			5718: Pixel = 99;
			5719: Pixel = 79;
			5720: Pixel = 78;
			5721: Pixel = 86;
			5722: Pixel = 93;
			5723: Pixel = 97;
			5724: Pixel = 99;
			5725: Pixel = 101;
			5726: Pixel = 101;
			5727: Pixel = 103;
			5728: Pixel = 100;
			5729: Pixel = 102;
			5730: Pixel = 107;
			5731: Pixel = 108;
			5732: Pixel = 110;
			5733: Pixel = 114;
			5734: Pixel = 109;
			5735: Pixel = 104;
			5736: Pixel = 198;
			5737: Pixel = 185;
			5738: Pixel = 123;
			5739: Pixel = 98;
			5740: Pixel = 100;
			5741: Pixel = 104;
			5742: Pixel = 99;
			5743: Pixel = 103;
			5744: Pixel = 118;
			5745: Pixel = 118;
			5746: Pixel = 123;
			5747: Pixel = 122;
			5748: Pixel = 116;
			5749: Pixel = 121;
			5750: Pixel = 120;
			5751: Pixel = 131;
			5752: Pixel = 133;
			5753: Pixel = 134;
			5754: Pixel = 128;
			5755: Pixel = 102;
			5756: Pixel = 129;
			5757: Pixel = 157;
			5758: Pixel = 172;
			5759: Pixel = 159;
			5760: Pixel = 154;
			5761: Pixel = 170;
			5762: Pixel = 164;
			5763: Pixel = 161;
			5764: Pixel = 175;
			5765: Pixel = 183;
			5766: Pixel = 179;
			5767: Pixel = 178;
			5768: Pixel = 179;
			5769: Pixel = 187;
			5770: Pixel = 184;
			5771: Pixel = 179;
			5772: Pixel = 184;
			5773: Pixel = 183;
			5774: Pixel = 169;
			5775: Pixel = 176;
			5776: Pixel = 191;
			5777: Pixel = 186;
			5778: Pixel = 192;
			5779: Pixel = 198;
			5780: Pixel = 196;
			5781: Pixel = 194;
			5782: Pixel = 197;
			5783: Pixel = 195;
			5784: Pixel = 195;
			5785: Pixel = 204;
			5786: Pixel = 194;
			5787: Pixel = 181;
			5788: Pixel = 190;
			5789: Pixel = 196;
			5790: Pixel = 198;
			5791: Pixel = 203;
			5792: Pixel = 202;
			5793: Pixel = 202;
			5794: Pixel = 205;
			5795: Pixel = 204;
			5796: Pixel = 209;
			5797: Pixel = 218;
			5798: Pixel = 181;
			5799: Pixel = 136;
			5800: Pixel = 148;
			5801: Pixel = 152;
			5802: Pixel = 154;
			5803: Pixel = 153;
			5804: Pixel = 150;
			5805: Pixel = 136;
			5806: Pixel = 95;
			5807: Pixel = 82;
			5808: Pixel = 156;
			5809: Pixel = 215;
			5810: Pixel = 195;
			5811: Pixel = 177;
			5812: Pixel = 205;
			5813: Pixel = 217;
			5814: Pixel = 209;
			5815: Pixel = 208;
			5816: Pixel = 202;
			5817: Pixel = 199;
			5818: Pixel = 203;
			5819: Pixel = 212;
			5820: Pixel = 217;
			5821: Pixel = 237;
			5822: Pixel = 148;
			5823: Pixel = 29;
			5824: Pixel = 49;
			5825: Pixel = 53;
			5826: Pixel = 57;
			5827: Pixel = 48;
			5828: Pixel = 46;
			5829: Pixel = 46;
			5830: Pixel = 45;
			5831: Pixel = 51;
			5832: Pixel = 54;
			5833: Pixel = 50;
			5834: Pixel = 33;
			5835: Pixel = 51;
			5836: Pixel = 124;
			5837: Pixel = 156;
			5838: Pixel = 146;
			5839: Pixel = 143;
			5840: Pixel = 157;
			5841: Pixel = 162;
			5842: Pixel = 159;
			5843: Pixel = 157;
			5844: Pixel = 157;
			5845: Pixel = 157;
			5846: Pixel = 157;
			5847: Pixel = 156;
			5848: Pixel = 154;
			5849: Pixel = 157;
			5850: Pixel = 99;
			5851: Pixel = 98;
			5852: Pixel = 99;
			5853: Pixel = 99;
			5854: Pixel = 99;
			5855: Pixel = 97;
			5856: Pixel = 93;
			5857: Pixel = 101;
			5858: Pixel = 126;
			5859: Pixel = 145;
			5860: Pixel = 158;
			5861: Pixel = 165;
			5862: Pixel = 167;
			5863: Pixel = 167;
			5864: Pixel = 168;
			5865: Pixel = 165;
			5866: Pixel = 152;
			5867: Pixel = 130;
			5868: Pixel = 100;
			5869: Pixel = 78;
			5870: Pixel = 79;
			5871: Pixel = 86;
			5872: Pixel = 93;
			5873: Pixel = 98;
			5874: Pixel = 99;
			5875: Pixel = 101;
			5876: Pixel = 102;
			5877: Pixel = 104;
			5878: Pixel = 101;
			5879: Pixel = 99;
			5880: Pixel = 107;
			5881: Pixel = 109;
			5882: Pixel = 111;
			5883: Pixel = 115;
			5884: Pixel = 105;
			5885: Pixel = 117;
			5886: Pixel = 213;
			5887: Pixel = 168;
			5888: Pixel = 114;
			5889: Pixel = 99;
			5890: Pixel = 94;
			5891: Pixel = 101;
			5892: Pixel = 109;
			5893: Pixel = 113;
			5894: Pixel = 112;
			5895: Pixel = 107;
			5896: Pixel = 117;
			5897: Pixel = 115;
			5898: Pixel = 119;
			5899: Pixel = 125;
			5900: Pixel = 129;
			5901: Pixel = 127;
			5902: Pixel = 120;
			5903: Pixel = 121;
			5904: Pixel = 105;
			5905: Pixel = 127;
			5906: Pixel = 161;
			5907: Pixel = 161;
			5908: Pixel = 149;
			5909: Pixel = 150;
			5910: Pixel = 155;
			5911: Pixel = 158;
			5912: Pixel = 164;
			5913: Pixel = 174;
			5914: Pixel = 172;
			5915: Pixel = 177;
			5916: Pixel = 181;
			5917: Pixel = 185;
			5918: Pixel = 174;
			5919: Pixel = 174;
			5920: Pixel = 183;
			5921: Pixel = 183;
			5922: Pixel = 174;
			5923: Pixel = 165;
			5924: Pixel = 180;
			5925: Pixel = 181;
			5926: Pixel = 189;
			5927: Pixel = 187;
			5928: Pixel = 185;
			5929: Pixel = 192;
			5930: Pixel = 195;
			5931: Pixel = 193;
			5932: Pixel = 196;
			5933: Pixel = 198;
			5934: Pixel = 200;
			5935: Pixel = 198;
			5936: Pixel = 170;
			5937: Pixel = 173;
			5938: Pixel = 196;
			5939: Pixel = 200;
			5940: Pixel = 202;
			5941: Pixel = 201;
			5942: Pixel = 201;
			5943: Pixel = 201;
			5944: Pixel = 198;
			5945: Pixel = 197;
			5946: Pixel = 202;
			5947: Pixel = 208;
			5948: Pixel = 221;
			5949: Pixel = 179;
			5950: Pixel = 144;
			5951: Pixel = 154;
			5952: Pixel = 151;
			5953: Pixel = 151;
			5954: Pixel = 139;
			5955: Pixel = 128;
			5956: Pixel = 146;
			5957: Pixel = 201;
			5958: Pixel = 212;
			5959: Pixel = 185;
			5960: Pixel = 187;
			5961: Pixel = 210;
			5962: Pixel = 214;
			5963: Pixel = 206;
			5964: Pixel = 204;
			5965: Pixel = 202;
			5966: Pixel = 199;
			5967: Pixel = 203;
			5968: Pixel = 207;
			5969: Pixel = 214;
			5970: Pixel = 217;
			5971: Pixel = 234;
			5972: Pixel = 129;
			5973: Pixel = 32;
			5974: Pixel = 50;
			5975: Pixel = 48;
			5976: Pixel = 53;
			5977: Pixel = 55;
			5978: Pixel = 49;
			5979: Pixel = 46;
			5980: Pixel = 49;
			5981: Pixel = 52;
			5982: Pixel = 55;
			5983: Pixel = 42;
			5984: Pixel = 31;
			5985: Pixel = 93;
			5986: Pixel = 152;
			5987: Pixel = 152;
			5988: Pixel = 144;
			5989: Pixel = 153;
			5990: Pixel = 161;
			5991: Pixel = 160;
			5992: Pixel = 158;
			5993: Pixel = 157;
			5994: Pixel = 155;
			5995: Pixel = 156;
			5996: Pixel = 155;
			5997: Pixel = 155;
			5998: Pixel = 154;
			5999: Pixel = 154;
			6000: Pixel = 100;
			6001: Pixel = 100;
			6002: Pixel = 101;
			6003: Pixel = 99;
			6004: Pixel = 100;
			6005: Pixel = 98;
			6006: Pixel = 97;
			6007: Pixel = 105;
			6008: Pixel = 128;
			6009: Pixel = 145;
			6010: Pixel = 155;
			6011: Pixel = 164;
			6012: Pixel = 167;
			6013: Pixel = 170;
			6014: Pixel = 168;
			6015: Pixel = 167;
			6016: Pixel = 153;
			6017: Pixel = 131;
			6018: Pixel = 103;
			6019: Pixel = 76;
			6020: Pixel = 79;
			6021: Pixel = 87;
			6022: Pixel = 92;
			6023: Pixel = 98;
			6024: Pixel = 100;
			6025: Pixel = 101;
			6026: Pixel = 101;
			6027: Pixel = 101;
			6028: Pixel = 100;
			6029: Pixel = 99;
			6030: Pixel = 103;
			6031: Pixel = 106;
			6032: Pixel = 109;
			6033: Pixel = 111;
			6034: Pixel = 96;
			6035: Pixel = 129;
			6036: Pixel = 212;
			6037: Pixel = 148;
			6038: Pixel = 122;
			6039: Pixel = 106;
			6040: Pixel = 99;
			6041: Pixel = 105;
			6042: Pixel = 105;
			6043: Pixel = 100;
			6044: Pixel = 102;
			6045: Pixel = 112;
			6046: Pixel = 115;
			6047: Pixel = 114;
			6048: Pixel = 125;
			6049: Pixel = 128;
			6050: Pixel = 119;
			6051: Pixel = 118;
			6052: Pixel = 118;
			6053: Pixel = 109;
			6054: Pixel = 129;
			6055: Pixel = 159;
			6056: Pixel = 158;
			6057: Pixel = 147;
			6058: Pixel = 148;
			6059: Pixel = 148;
			6060: Pixel = 146;
			6061: Pixel = 152;
			6062: Pixel = 171;
			6063: Pixel = 174;
			6064: Pixel = 178;
			6065: Pixel = 175;
			6066: Pixel = 170;
			6067: Pixel = 168;
			6068: Pixel = 180;
			6069: Pixel = 181;
			6070: Pixel = 177;
			6071: Pixel = 173;
			6072: Pixel = 167;
			6073: Pixel = 177;
			6074: Pixel = 186;
			6075: Pixel = 182;
			6076: Pixel = 181;
			6077: Pixel = 183;
			6078: Pixel = 186;
			6079: Pixel = 183;
			6080: Pixel = 187;
			6081: Pixel = 192;
			6082: Pixel = 197;
			6083: Pixel = 204;
			6084: Pixel = 193;
			6085: Pixel = 173;
			6086: Pixel = 178;
			6087: Pixel = 193;
			6088: Pixel = 193;
			6089: Pixel = 197;
			6090: Pixel = 197;
			6091: Pixel = 197;
			6092: Pixel = 200;
			6093: Pixel = 198;
			6094: Pixel = 199;
			6095: Pixel = 195;
			6096: Pixel = 194;
			6097: Pixel = 197;
			6098: Pixel = 203;
			6099: Pixel = 206;
			6100: Pixel = 155;
			6101: Pixel = 153;
			6102: Pixel = 147;
			6103: Pixel = 141;
			6104: Pixel = 158;
			6105: Pixel = 196;
			6106: Pixel = 211;
			6107: Pixel = 195;
			6108: Pixel = 182;
			6109: Pixel = 196;
			6110: Pixel = 211;
			6111: Pixel = 209;
			6112: Pixel = 204;
			6113: Pixel = 201;
			6114: Pixel = 201;
			6115: Pixel = 201;
			6116: Pixel = 202;
			6117: Pixel = 206;
			6118: Pixel = 212;
			6119: Pixel = 215;
			6120: Pixel = 218;
			6121: Pixel = 229;
			6122: Pixel = 98;
			6123: Pixel = 33;
			6124: Pixel = 54;
			6125: Pixel = 49;
			6126: Pixel = 48;
			6127: Pixel = 52;
			6128: Pixel = 47;
			6129: Pixel = 42;
			6130: Pixel = 46;
			6131: Pixel = 52;
			6132: Pixel = 50;
			6133: Pixel = 41;
			6134: Pixel = 65;
			6135: Pixel = 134;
			6136: Pixel = 155;
			6137: Pixel = 147;
			6138: Pixel = 147;
			6139: Pixel = 159;
			6140: Pixel = 160;
			6141: Pixel = 159;
			6142: Pixel = 157;
			6143: Pixel = 157;
			6144: Pixel = 156;
			6145: Pixel = 156;
			6146: Pixel = 156;
			6147: Pixel = 155;
			6148: Pixel = 153;
			6149: Pixel = 154;
			6150: Pixel = 100;
			6151: Pixel = 99;
			6152: Pixel = 98;
			6153: Pixel = 99;
			6154: Pixel = 100;
			6155: Pixel = 98;
			6156: Pixel = 97;
			6157: Pixel = 108;
			6158: Pixel = 129;
			6159: Pixel = 147;
			6160: Pixel = 158;
			6161: Pixel = 165;
			6162: Pixel = 169;
			6163: Pixel = 171;
			6164: Pixel = 172;
			6165: Pixel = 169;
			6166: Pixel = 154;
			6167: Pixel = 132;
			6168: Pixel = 100;
			6169: Pixel = 77;
			6170: Pixel = 79;
			6171: Pixel = 90;
			6172: Pixel = 94;
			6173: Pixel = 98;
			6174: Pixel = 98;
			6175: Pixel = 101;
			6176: Pixel = 101;
			6177: Pixel = 101;
			6178: Pixel = 99;
			6179: Pixel = 100;
			6180: Pixel = 102;
			6181: Pixel = 107;
			6182: Pixel = 107;
			6183: Pixel = 108;
			6184: Pixel = 89;
			6185: Pixel = 151;
			6186: Pixel = 208;
			6187: Pixel = 148;
			6188: Pixel = 128;
			6189: Pixel = 108;
			6190: Pixel = 105;
			6191: Pixel = 105;
			6192: Pixel = 104;
			6193: Pixel = 101;
			6194: Pixel = 104;
			6195: Pixel = 110;
			6196: Pixel = 107;
			6197: Pixel = 118;
			6198: Pixel = 121;
			6199: Pixel = 115;
			6200: Pixel = 118;
			6201: Pixel = 121;
			6202: Pixel = 113;
			6203: Pixel = 141;
			6204: Pixel = 150;
			6205: Pixel = 148;
			6206: Pixel = 146;
			6207: Pixel = 147;
			6208: Pixel = 148;
			6209: Pixel = 138;
			6210: Pixel = 154;
			6211: Pixel = 165;
			6212: Pixel = 161;
			6213: Pixel = 176;
			6214: Pixel = 174;
			6215: Pixel = 165;
			6216: Pixel = 165;
			6217: Pixel = 169;
			6218: Pixel = 178;
			6219: Pixel = 184;
			6220: Pixel = 159;
			6221: Pixel = 164;
			6222: Pixel = 182;
			6223: Pixel = 174;
			6224: Pixel = 174;
			6225: Pixel = 183;
			6226: Pixel = 178;
			6227: Pixel = 177;
			6228: Pixel = 175;
			6229: Pixel = 178;
			6230: Pixel = 183;
			6231: Pixel = 191;
			6232: Pixel = 178;
			6233: Pixel = 180;
			6234: Pixel = 175;
			6235: Pixel = 185;
			6236: Pixel = 188;
			6237: Pixel = 183;
			6238: Pixel = 186;
			6239: Pixel = 192;
			6240: Pixel = 194;
			6241: Pixel = 196;
			6242: Pixel = 191;
			6243: Pixel = 191;
			6244: Pixel = 192;
			6245: Pixel = 195;
			6246: Pixel = 188;
			6247: Pixel = 188;
			6248: Pixel = 189;
			6249: Pixel = 203;
			6250: Pixel = 169;
			6251: Pixel = 141;
			6252: Pixel = 156;
			6253: Pixel = 180;
			6254: Pixel = 205;
			6255: Pixel = 201;
			6256: Pixel = 185;
			6257: Pixel = 187;
			6258: Pixel = 206;
			6259: Pixel = 210;
			6260: Pixel = 204;
			6261: Pixel = 201;
			6262: Pixel = 200;
			6263: Pixel = 200;
			6264: Pixel = 202;
			6265: Pixel = 204;
			6266: Pixel = 204;
			6267: Pixel = 206;
			6268: Pixel = 210;
			6269: Pixel = 216;
			6270: Pixel = 222;
			6271: Pixel = 218;
			6272: Pixel = 74;
			6273: Pixel = 42;
			6274: Pixel = 55;
			6275: Pixel = 53;
			6276: Pixel = 50;
			6277: Pixel = 48;
			6278: Pixel = 42;
			6279: Pixel = 44;
			6280: Pixel = 49;
			6281: Pixel = 51;
			6282: Pixel = 55;
			6283: Pixel = 61;
			6284: Pixel = 109;
			6285: Pixel = 151;
			6286: Pixel = 148;
			6287: Pixel = 145;
			6288: Pixel = 154;
			6289: Pixel = 160;
			6290: Pixel = 160;
			6291: Pixel = 159;
			6292: Pixel = 158;
			6293: Pixel = 157;
			6294: Pixel = 158;
			6295: Pixel = 156;
			6296: Pixel = 154;
			6297: Pixel = 154;
			6298: Pixel = 154;
			6299: Pixel = 152;
			6300: Pixel = 100;
			6301: Pixel = 100;
			6302: Pixel = 101;
			6303: Pixel = 98;
			6304: Pixel = 100;
			6305: Pixel = 100;
			6306: Pixel = 97;
			6307: Pixel = 108;
			6308: Pixel = 128;
			6309: Pixel = 148;
			6310: Pixel = 161;
			6311: Pixel = 167;
			6312: Pixel = 171;
			6313: Pixel = 172;
			6314: Pixel = 173;
			6315: Pixel = 171;
			6316: Pixel = 156;
			6317: Pixel = 132;
			6318: Pixel = 101;
			6319: Pixel = 78;
			6320: Pixel = 79;
			6321: Pixel = 91;
			6322: Pixel = 92;
			6323: Pixel = 97;
			6324: Pixel = 99;
			6325: Pixel = 100;
			6326: Pixel = 99;
			6327: Pixel = 98;
			6328: Pixel = 97;
			6329: Pixel = 100;
			6330: Pixel = 101;
			6331: Pixel = 104;
			6332: Pixel = 106;
			6333: Pixel = 104;
			6334: Pixel = 86;
			6335: Pixel = 175;
			6336: Pixel = 205;
			6337: Pixel = 156;
			6338: Pixel = 131;
			6339: Pixel = 111;
			6340: Pixel = 100;
			6341: Pixel = 106;
			6342: Pixel = 107;
			6343: Pixel = 106;
			6344: Pixel = 108;
			6345: Pixel = 111;
			6346: Pixel = 114;
			6347: Pixel = 119;
			6348: Pixel = 113;
			6349: Pixel = 123;
			6350: Pixel = 126;
			6351: Pixel = 112;
			6352: Pixel = 134;
			6353: Pixel = 152;
			6354: Pixel = 153;
			6355: Pixel = 139;
			6356: Pixel = 144;
			6357: Pixel = 144;
			6358: Pixel = 132;
			6359: Pixel = 152;
			6360: Pixel = 159;
			6361: Pixel = 162;
			6362: Pixel = 166;
			6363: Pixel = 156;
			6364: Pixel = 164;
			6365: Pixel = 174;
			6366: Pixel = 172;
			6367: Pixel = 175;
			6368: Pixel = 164;
			6369: Pixel = 157;
			6370: Pixel = 169;
			6371: Pixel = 176;
			6372: Pixel = 173;
			6373: Pixel = 179;
			6374: Pixel = 175;
			6375: Pixel = 174;
			6376: Pixel = 174;
			6377: Pixel = 179;
			6378: Pixel = 179;
			6379: Pixel = 187;
			6380: Pixel = 189;
			6381: Pixel = 176;
			6382: Pixel = 170;
			6383: Pixel = 180;
			6384: Pixel = 189;
			6385: Pixel = 183;
			6386: Pixel = 178;
			6387: Pixel = 190;
			6388: Pixel = 190;
			6389: Pixel = 194;
			6390: Pixel = 192;
			6391: Pixel = 192;
			6392: Pixel = 183;
			6393: Pixel = 187;
			6394: Pixel = 188;
			6395: Pixel = 187;
			6396: Pixel = 185;
			6397: Pixel = 184;
			6398: Pixel = 187;
			6399: Pixel = 188;
			6400: Pixel = 189;
			6401: Pixel = 171;
			6402: Pixel = 202;
			6403: Pixel = 201;
			6404: Pixel = 186;
			6405: Pixel = 190;
			6406: Pixel = 201;
			6407: Pixel = 207;
			6408: Pixel = 208;
			6409: Pixel = 202;
			6410: Pixel = 200;
			6411: Pixel = 199;
			6412: Pixel = 200;
			6413: Pixel = 203;
			6414: Pixel = 205;
			6415: Pixel = 204;
			6416: Pixel = 200;
			6417: Pixel = 201;
			6418: Pixel = 210;
			6419: Pixel = 215;
			6420: Pixel = 227;
			6421: Pixel = 203;
			6422: Pixel = 52;
			6423: Pixel = 44;
			6424: Pixel = 51;
			6425: Pixel = 51;
			6426: Pixel = 55;
			6427: Pixel = 48;
			6428: Pixel = 43;
			6429: Pixel = 48;
			6430: Pixel = 49;
			6431: Pixel = 55;
			6432: Pixel = 63;
			6433: Pixel = 89;
			6434: Pixel = 139;
			6435: Pixel = 151;
			6436: Pixel = 143;
			6437: Pixel = 150;
			6438: Pixel = 159;
			6439: Pixel = 161;
			6440: Pixel = 159;
			6441: Pixel = 159;
			6442: Pixel = 157;
			6443: Pixel = 156;
			6444: Pixel = 157;
			6445: Pixel = 155;
			6446: Pixel = 154;
			6447: Pixel = 155;
			6448: Pixel = 153;
			6449: Pixel = 154;
			6450: Pixel = 100;
			6451: Pixel = 99;
			6452: Pixel = 99;
			6453: Pixel = 96;
			6454: Pixel = 99;
			6455: Pixel = 99;
			6456: Pixel = 100;
			6457: Pixel = 108;
			6458: Pixel = 127;
			6459: Pixel = 147;
			6460: Pixel = 161;
			6461: Pixel = 169;
			6462: Pixel = 172;
			6463: Pixel = 174;
			6464: Pixel = 173;
			6465: Pixel = 170;
			6466: Pixel = 156;
			6467: Pixel = 132;
			6468: Pixel = 102;
			6469: Pixel = 77;
			6470: Pixel = 77;
			6471: Pixel = 85;
			6472: Pixel = 92;
			6473: Pixel = 95;
			6474: Pixel = 98;
			6475: Pixel = 100;
			6476: Pixel = 99;
			6477: Pixel = 98;
			6478: Pixel = 98;
			6479: Pixel = 98;
			6480: Pixel = 98;
			6481: Pixel = 104;
			6482: Pixel = 105;
			6483: Pixel = 99;
			6484: Pixel = 92;
			6485: Pixel = 195;
			6486: Pixel = 200;
			6487: Pixel = 161;
			6488: Pixel = 139;
			6489: Pixel = 119;
			6490: Pixel = 112;
			6491: Pixel = 109;
			6492: Pixel = 102;
			6493: Pixel = 105;
			6494: Pixel = 110;
			6495: Pixel = 115;
			6496: Pixel = 116;
			6497: Pixel = 120;
			6498: Pixel = 123;
			6499: Pixel = 127;
			6500: Pixel = 106;
			6501: Pixel = 132;
			6502: Pixel = 152;
			6503: Pixel = 144;
			6504: Pixel = 141;
			6505: Pixel = 149;
			6506: Pixel = 134;
			6507: Pixel = 130;
			6508: Pixel = 147;
			6509: Pixel = 149;
			6510: Pixel = 157;
			6511: Pixel = 160;
			6512: Pixel = 151;
			6513: Pixel = 162;
			6514: Pixel = 166;
			6515: Pixel = 174;
			6516: Pixel = 180;
			6517: Pixel = 160;
			6518: Pixel = 156;
			6519: Pixel = 173;
			6520: Pixel = 179;
			6521: Pixel = 170;
			6522: Pixel = 172;
			6523: Pixel = 173;
			6524: Pixel = 175;
			6525: Pixel = 174;
			6526: Pixel = 169;
			6527: Pixel = 172;
			6528: Pixel = 182;
			6529: Pixel = 186;
			6530: Pixel = 180;
			6531: Pixel = 181;
			6532: Pixel = 183;
			6533: Pixel = 181;
			6534: Pixel = 182;
			6535: Pixel = 189;
			6536: Pixel = 189;
			6537: Pixel = 188;
			6538: Pixel = 191;
			6539: Pixel = 187;
			6540: Pixel = 183;
			6541: Pixel = 177;
			6542: Pixel = 180;
			6543: Pixel = 186;
			6544: Pixel = 183;
			6545: Pixel = 182;
			6546: Pixel = 183;
			6547: Pixel = 170;
			6548: Pixel = 175;
			6549: Pixel = 187;
			6550: Pixel = 197;
			6551: Pixel = 195;
			6552: Pixel = 193;
			6553: Pixel = 191;
			6554: Pixel = 198;
			6555: Pixel = 208;
			6556: Pixel = 207;
			6557: Pixel = 199;
			6558: Pixel = 201;
			6559: Pixel = 200;
			6560: Pixel = 199;
			6561: Pixel = 197;
			6562: Pixel = 201;
			6563: Pixel = 203;
			6564: Pixel = 205;
			6565: Pixel = 202;
			6566: Pixel = 190;
			6567: Pixel = 203;
			6568: Pixel = 209;
			6569: Pixel = 213;
			6570: Pixel = 230;
			6571: Pixel = 170;
			6572: Pixel = 32;
			6573: Pixel = 45;
			6574: Pixel = 46;
			6575: Pixel = 48;
			6576: Pixel = 51;
			6577: Pixel = 45;
			6578: Pixel = 44;
			6579: Pixel = 51;
			6580: Pixel = 53;
			6581: Pixel = 54;
			6582: Pixel = 74;
			6583: Pixel = 124;
			6584: Pixel = 153;
			6585: Pixel = 147;
			6586: Pixel = 145;
			6587: Pixel = 156;
			6588: Pixel = 161;
			6589: Pixel = 160;
			6590: Pixel = 159;
			6591: Pixel = 158;
			6592: Pixel = 157;
			6593: Pixel = 156;
			6594: Pixel = 157;
			6595: Pixel = 156;
			6596: Pixel = 156;
			6597: Pixel = 155;
			6598: Pixel = 155;
			6599: Pixel = 156;
			6600: Pixel = 99;
			6601: Pixel = 96;
			6602: Pixel = 99;
			6603: Pixel = 97;
			6604: Pixel = 96;
			6605: Pixel = 97;
			6606: Pixel = 97;
			6607: Pixel = 104;
			6608: Pixel = 126;
			6609: Pixel = 146;
			6610: Pixel = 160;
			6611: Pixel = 170;
			6612: Pixel = 173;
			6613: Pixel = 173;
			6614: Pixel = 173;
			6615: Pixel = 170;
			6616: Pixel = 154;
			6617: Pixel = 132;
			6618: Pixel = 103;
			6619: Pixel = 77;
			6620: Pixel = 78;
			6621: Pixel = 87;
			6622: Pixel = 93;
			6623: Pixel = 97;
			6624: Pixel = 98;
			6625: Pixel = 97;
			6626: Pixel = 98;
			6627: Pixel = 99;
			6628: Pixel = 98;
			6629: Pixel = 98;
			6630: Pixel = 101;
			6631: Pixel = 104;
			6632: Pixel = 105;
			6633: Pixel = 99;
			6634: Pixel = 97;
			6635: Pixel = 201;
			6636: Pixel = 195;
			6637: Pixel = 160;
			6638: Pixel = 141;
			6639: Pixel = 131;
			6640: Pixel = 124;
			6641: Pixel = 115;
			6642: Pixel = 105;
			6643: Pixel = 106;
			6644: Pixel = 110;
			6645: Pixel = 103;
			6646: Pixel = 112;
			6647: Pixel = 121;
			6648: Pixel = 119;
			6649: Pixel = 112;
			6650: Pixel = 129;
			6651: Pixel = 145;
			6652: Pixel = 147;
			6653: Pixel = 137;
			6654: Pixel = 145;
			6655: Pixel = 135;
			6656: Pixel = 130;
			6657: Pixel = 152;
			6658: Pixel = 149;
			6659: Pixel = 155;
			6660: Pixel = 141;
			6661: Pixel = 141;
			6662: Pixel = 155;
			6663: Pixel = 170;
			6664: Pixel = 178;
			6665: Pixel = 166;
			6666: Pixel = 149;
			6667: Pixel = 164;
			6668: Pixel = 179;
			6669: Pixel = 169;
			6670: Pixel = 166;
			6671: Pixel = 173;
			6672: Pixel = 176;
			6673: Pixel = 176;
			6674: Pixel = 171;
			6675: Pixel = 176;
			6676: Pixel = 173;
			6677: Pixel = 168;
			6678: Pixel = 170;
			6679: Pixel = 174;
			6680: Pixel = 184;
			6681: Pixel = 182;
			6682: Pixel = 177;
			6683: Pixel = 182;
			6684: Pixel = 176;
			6685: Pixel = 183;
			6686: Pixel = 192;
			6687: Pixel = 187;
			6688: Pixel = 183;
			6689: Pixel = 182;
			6690: Pixel = 179;
			6691: Pixel = 172;
			6692: Pixel = 174;
			6693: Pixel = 184;
			6694: Pixel = 181;
			6695: Pixel = 172;
			6696: Pixel = 162;
			6697: Pixel = 166;
			6698: Pixel = 190;
			6699: Pixel = 193;
			6700: Pixel = 181;
			6701: Pixel = 184;
			6702: Pixel = 196;
			6703: Pixel = 203;
			6704: Pixel = 208;
			6705: Pixel = 207;
			6706: Pixel = 197;
			6707: Pixel = 196;
			6708: Pixel = 200;
			6709: Pixel = 199;
			6710: Pixel = 197;
			6711: Pixel = 201;
			6712: Pixel = 203;
			6713: Pixel = 204;
			6714: Pixel = 206;
			6715: Pixel = 179;
			6716: Pixel = 173;
			6717: Pixel = 198;
			6718: Pixel = 208;
			6719: Pixel = 209;
			6720: Pixel = 227;
			6721: Pixel = 120;
			6722: Pixel = 28;
			6723: Pixel = 45;
			6724: Pixel = 46;
			6725: Pixel = 49;
			6726: Pixel = 56;
			6727: Pixel = 46;
			6728: Pixel = 46;
			6729: Pixel = 55;
			6730: Pixel = 51;
			6731: Pixel = 42;
			6732: Pixel = 97;
			6733: Pixel = 149;
			6734: Pixel = 150;
			6735: Pixel = 144;
			6736: Pixel = 152;
			6737: Pixel = 159;
			6738: Pixel = 160;
			6739: Pixel = 160;
			6740: Pixel = 159;
			6741: Pixel = 160;
			6742: Pixel = 158;
			6743: Pixel = 157;
			6744: Pixel = 158;
			6745: Pixel = 158;
			6746: Pixel = 157;
			6747: Pixel = 156;
			6748: Pixel = 157;
			6749: Pixel = 157;
			6750: Pixel = 97;
			6751: Pixel = 99;
			6752: Pixel = 98;
			6753: Pixel = 97;
			6754: Pixel = 98;
			6755: Pixel = 98;
			6756: Pixel = 95;
			6757: Pixel = 105;
			6758: Pixel = 127;
			6759: Pixel = 147;
			6760: Pixel = 161;
			6761: Pixel = 170;
			6762: Pixel = 172;
			6763: Pixel = 173;
			6764: Pixel = 173;
			6765: Pixel = 170;
			6766: Pixel = 154;
			6767: Pixel = 134;
			6768: Pixel = 103;
			6769: Pixel = 79;
			6770: Pixel = 81;
			6771: Pixel = 90;
			6772: Pixel = 94;
			6773: Pixel = 95;
			6774: Pixel = 100;
			6775: Pixel = 101;
			6776: Pixel = 97;
			6777: Pixel = 99;
			6778: Pixel = 98;
			6779: Pixel = 98;
			6780: Pixel = 100;
			6781: Pixel = 102;
			6782: Pixel = 104;
			6783: Pixel = 97;
			6784: Pixel = 100;
			6785: Pixel = 204;
			6786: Pixel = 190;
			6787: Pixel = 166;
			6788: Pixel = 151;
			6789: Pixel = 139;
			6790: Pixel = 133;
			6791: Pixel = 117;
			6792: Pixel = 108;
			6793: Pixel = 101;
			6794: Pixel = 105;
			6795: Pixel = 109;
			6796: Pixel = 121;
			6797: Pixel = 114;
			6798: Pixel = 100;
			6799: Pixel = 134;
			6800: Pixel = 143;
			6801: Pixel = 140;
			6802: Pixel = 142;
			6803: Pixel = 145;
			6804: Pixel = 127;
			6805: Pixel = 125;
			6806: Pixel = 148;
			6807: Pixel = 148;
			6808: Pixel = 154;
			6809: Pixel = 148;
			6810: Pixel = 139;
			6811: Pixel = 151;
			6812: Pixel = 149;
			6813: Pixel = 159;
			6814: Pixel = 161;
			6815: Pixel = 154;
			6816: Pixel = 161;
			6817: Pixel = 174;
			6818: Pixel = 173;
			6819: Pixel = 169;
			6820: Pixel = 163;
			6821: Pixel = 168;
			6822: Pixel = 175;
			6823: Pixel = 175;
			6824: Pixel = 170;
			6825: Pixel = 162;
			6826: Pixel = 165;
			6827: Pixel = 170;
			6828: Pixel = 168;
			6829: Pixel = 172;
			6830: Pixel = 171;
			6831: Pixel = 169;
			6832: Pixel = 176;
			6833: Pixel = 183;
			6834: Pixel = 185;
			6835: Pixel = 179;
			6836: Pixel = 186;
			6837: Pixel = 183;
			6838: Pixel = 175;
			6839: Pixel = 176;
			6840: Pixel = 183;
			6841: Pixel = 181;
			6842: Pixel = 172;
			6843: Pixel = 172;
			6844: Pixel = 171;
			6845: Pixel = 160;
			6846: Pixel = 180;
			6847: Pixel = 197;
			6848: Pixel = 189;
			6849: Pixel = 184;
			6850: Pixel = 191;
			6851: Pixel = 202;
			6852: Pixel = 205;
			6853: Pixel = 202;
			6854: Pixel = 200;
			6855: Pixel = 197;
			6856: Pixel = 196;
			6857: Pixel = 199;
			6858: Pixel = 199;
			6859: Pixel = 199;
			6860: Pixel = 200;
			6861: Pixel = 202;
			6862: Pixel = 204;
			6863: Pixel = 206;
			6864: Pixel = 188;
			6865: Pixel = 156;
			6866: Pixel = 163;
			6867: Pixel = 188;
			6868: Pixel = 183;
			6869: Pixel = 205;
			6870: Pixel = 206;
			6871: Pixel = 64;
			6872: Pixel = 40;
			6873: Pixel = 48;
			6874: Pixel = 47;
			6875: Pixel = 51;
			6876: Pixel = 50;
			6877: Pixel = 44;
			6878: Pixel = 47;
			6879: Pixel = 48;
			6880: Pixel = 53;
			6881: Pixel = 65;
			6882: Pixel = 128;
			6883: Pixel = 155;
			6884: Pixel = 146;
			6885: Pixel = 149;
			6886: Pixel = 159;
			6887: Pixel = 160;
			6888: Pixel = 161;
			6889: Pixel = 160;
			6890: Pixel = 159;
			6891: Pixel = 160;
			6892: Pixel = 157;
			6893: Pixel = 157;
			6894: Pixel = 157;
			6895: Pixel = 156;
			6896: Pixel = 158;
			6897: Pixel = 158;
			6898: Pixel = 156;
			6899: Pixel = 156;
			6900: Pixel = 97;
			6901: Pixel = 96;
			6902: Pixel = 95;
			6903: Pixel = 94;
			6904: Pixel = 96;
			6905: Pixel = 96;
			6906: Pixel = 97;
			6907: Pixel = 104;
			6908: Pixel = 129;
			6909: Pixel = 151;
			6910: Pixel = 163;
			6911: Pixel = 171;
			6912: Pixel = 171;
			6913: Pixel = 171;
			6914: Pixel = 170;
			6915: Pixel = 168;
			6916: Pixel = 155;
			6917: Pixel = 133;
			6918: Pixel = 101;
			6919: Pixel = 79;
			6920: Pixel = 79;
			6921: Pixel = 90;
			6922: Pixel = 95;
			6923: Pixel = 98;
			6924: Pixel = 100;
			6925: Pixel = 98;
			6926: Pixel = 99;
			6927: Pixel = 99;
			6928: Pixel = 98;
			6929: Pixel = 98;
			6930: Pixel = 100;
			6931: Pixel = 102;
			6932: Pixel = 102;
			6933: Pixel = 95;
			6934: Pixel = 100;
			6935: Pixel = 201;
			6936: Pixel = 188;
			6937: Pixel = 165;
			6938: Pixel = 158;
			6939: Pixel = 145;
			6940: Pixel = 138;
			6941: Pixel = 130;
			6942: Pixel = 114;
			6943: Pixel = 95;
			6944: Pixel = 95;
			6945: Pixel = 111;
			6946: Pixel = 114;
			6947: Pixel = 106;
			6948: Pixel = 129;
			6949: Pixel = 143;
			6950: Pixel = 138;
			6951: Pixel = 133;
			6952: Pixel = 146;
			6953: Pixel = 125;
			6954: Pixel = 119;
			6955: Pixel = 146;
			6956: Pixel = 152;
			6957: Pixel = 147;
			6958: Pixel = 142;
			6959: Pixel = 148;
			6960: Pixel = 153;
			6961: Pixel = 150;
			6962: Pixel = 146;
			6963: Pixel = 149;
			6964: Pixel = 147;
			6965: Pixel = 157;
			6966: Pixel = 176;
			6967: Pixel = 169;
			6968: Pixel = 163;
			6969: Pixel = 166;
			6970: Pixel = 171;
			6971: Pixel = 166;
			6972: Pixel = 162;
			6973: Pixel = 168;
			6974: Pixel = 163;
			6975: Pixel = 166;
			6976: Pixel = 166;
			6977: Pixel = 163;
			6978: Pixel = 162;
			6979: Pixel = 157;
			6980: Pixel = 168;
			6981: Pixel = 174;
			6982: Pixel = 174;
			6983: Pixel = 172;
			6984: Pixel = 183;
			6985: Pixel = 183;
			6986: Pixel = 173;
			6987: Pixel = 175;
			6988: Pixel = 174;
			6989: Pixel = 168;
			6990: Pixel = 178;
			6991: Pixel = 181;
			6992: Pixel = 161;
			6993: Pixel = 153;
			6994: Pixel = 173;
			6995: Pixel = 189;
			6996: Pixel = 190;
			6997: Pixel = 183;
			6998: Pixel = 190;
			6999: Pixel = 201;
			7000: Pixel = 205;
			7001: Pixel = 200;
			7002: Pixel = 196;
			7003: Pixel = 192;
			7004: Pixel = 190;
			7005: Pixel = 194;
			7006: Pixel = 197;
			7007: Pixel = 200;
			7008: Pixel = 200;
			7009: Pixel = 199;
			7010: Pixel = 201;
			7011: Pixel = 204;
			7012: Pixel = 206;
			7013: Pixel = 201;
			7014: Pixel = 159;
			7015: Pixel = 158;
			7016: Pixel = 178;
			7017: Pixel = 143;
			7018: Pixel = 159;
			7019: Pixel = 208;
			7020: Pixel = 155;
			7021: Pixel = 32;
			7022: Pixel = 48;
			7023: Pixel = 55;
			7024: Pixel = 53;
			7025: Pixel = 49;
			7026: Pixel = 43;
			7027: Pixel = 47;
			7028: Pixel = 46;
			7029: Pixel = 48;
			7030: Pixel = 72;
			7031: Pixel = 109;
			7032: Pixel = 149;
			7033: Pixel = 148;
			7034: Pixel = 144;
			7035: Pixel = 155;
			7036: Pixel = 159;
			7037: Pixel = 160;
			7038: Pixel = 159;
			7039: Pixel = 158;
			7040: Pixel = 159;
			7041: Pixel = 159;
			7042: Pixel = 157;
			7043: Pixel = 157;
			7044: Pixel = 157;
			7045: Pixel = 157;
			7046: Pixel = 158;
			7047: Pixel = 158;
			7048: Pixel = 156;
			7049: Pixel = 157;
			7050: Pixel = 98;
			7051: Pixel = 95;
			7052: Pixel = 93;
			7053: Pixel = 95;
			7054: Pixel = 94;
			7055: Pixel = 95;
			7056: Pixel = 96;
			7057: Pixel = 106;
			7058: Pixel = 130;
			7059: Pixel = 150;
			7060: Pixel = 162;
			7061: Pixel = 169;
			7062: Pixel = 171;
			7063: Pixel = 171;
			7064: Pixel = 171;
			7065: Pixel = 167;
			7066: Pixel = 156;
			7067: Pixel = 135;
			7068: Pixel = 102;
			7069: Pixel = 78;
			7070: Pixel = 78;
			7071: Pixel = 88;
			7072: Pixel = 95;
			7073: Pixel = 97;
			7074: Pixel = 99;
			7075: Pixel = 99;
			7076: Pixel = 97;
			7077: Pixel = 97;
			7078: Pixel = 98;
			7079: Pixel = 98;
			7080: Pixel = 101;
			7081: Pixel = 100;
			7082: Pixel = 100;
			7083: Pixel = 89;
			7084: Pixel = 106;
			7085: Pixel = 203;
			7086: Pixel = 182;
			7087: Pixel = 166;
			7088: Pixel = 157;
			7089: Pixel = 147;
			7090: Pixel = 137;
			7091: Pixel = 135;
			7092: Pixel = 109;
			7093: Pixel = 100;
			7094: Pixel = 102;
			7095: Pixel = 108;
			7096: Pixel = 101;
			7097: Pixel = 131;
			7098: Pixel = 145;
			7099: Pixel = 132;
			7100: Pixel = 133;
			7101: Pixel = 140;
			7102: Pixel = 121;
			7103: Pixel = 120;
			7104: Pixel = 143;
			7105: Pixel = 141;
			7106: Pixel = 146;
			7107: Pixel = 141;
			7108: Pixel = 141;
			7109: Pixel = 142;
			7110: Pixel = 143;
			7111: Pixel = 155;
			7112: Pixel = 153;
			7113: Pixel = 140;
			7114: Pixel = 160;
			7115: Pixel = 163;
			7116: Pixel = 154;
			7117: Pixel = 159;
			7118: Pixel = 171;
			7119: Pixel = 167;
			7120: Pixel = 163;
			7121: Pixel = 163;
			7122: Pixel = 160;
			7123: Pixel = 161;
			7124: Pixel = 170;
			7125: Pixel = 159;
			7126: Pixel = 157;
			7127: Pixel = 160;
			7128: Pixel = 161;
			7129: Pixel = 166;
			7130: Pixel = 167;
			7131: Pixel = 171;
			7132: Pixel = 172;
			7133: Pixel = 165;
			7134: Pixel = 171;
			7135: Pixel = 176;
			7136: Pixel = 172;
			7137: Pixel = 168;
			7138: Pixel = 172;
			7139: Pixel = 166;
			7140: Pixel = 166;
			7141: Pixel = 162;
			7142: Pixel = 163;
			7143: Pixel = 182;
			7144: Pixel = 187;
			7145: Pixel = 179;
			7146: Pixel = 185;
			7147: Pixel = 197;
			7148: Pixel = 207;
			7149: Pixel = 204;
			7150: Pixel = 197;
			7151: Pixel = 192;
			7152: Pixel = 191;
			7153: Pixel = 193;
			7154: Pixel = 192;
			7155: Pixel = 197;
			7156: Pixel = 199;
			7157: Pixel = 201;
			7158: Pixel = 200;
			7159: Pixel = 201;
			7160: Pixel = 203;
			7161: Pixel = 206;
			7162: Pixel = 211;
			7163: Pixel = 173;
			7164: Pixel = 156;
			7165: Pixel = 177;
			7166: Pixel = 145;
			7167: Pixel = 145;
			7168: Pixel = 172;
			7169: Pixel = 211;
			7170: Pixel = 101;
			7171: Pixel = 27;
			7172: Pixel = 43;
			7173: Pixel = 51;
			7174: Pixel = 55;
			7175: Pixel = 42;
			7176: Pixel = 44;
			7177: Pixel = 52;
			7178: Pixel = 46;
			7179: Pixel = 58;
			7180: Pixel = 88;
			7181: Pixel = 141;
			7182: Pixel = 154;
			7183: Pixel = 144;
			7184: Pixel = 149;
			7185: Pixel = 159;
			7186: Pixel = 160;
			7187: Pixel = 161;
			7188: Pixel = 160;
			7189: Pixel = 157;
			7190: Pixel = 157;
			7191: Pixel = 158;
			7192: Pixel = 159;
			7193: Pixel = 158;
			7194: Pixel = 156;
			7195: Pixel = 156;
			7196: Pixel = 157;
			7197: Pixel = 157;
			7198: Pixel = 156;
			7199: Pixel = 157;
			7200: Pixel = 97;
			7201: Pixel = 97;
			7202: Pixel = 92;
			7203: Pixel = 96;
			7204: Pixel = 94;
			7205: Pixel = 94;
			7206: Pixel = 96;
			7207: Pixel = 108;
			7208: Pixel = 131;
			7209: Pixel = 149;
			7210: Pixel = 163;
			7211: Pixel = 169;
			7212: Pixel = 171;
			7213: Pixel = 170;
			7214: Pixel = 171;
			7215: Pixel = 169;
			7216: Pixel = 156;
			7217: Pixel = 136;
			7218: Pixel = 104;
			7219: Pixel = 79;
			7220: Pixel = 80;
			7221: Pixel = 90;
			7222: Pixel = 94;
			7223: Pixel = 98;
			7224: Pixel = 98;
			7225: Pixel = 97;
			7226: Pixel = 98;
			7227: Pixel = 98;
			7228: Pixel = 97;
			7229: Pixel = 100;
			7230: Pixel = 99;
			7231: Pixel = 99;
			7232: Pixel = 100;
			7233: Pixel = 83;
			7234: Pixel = 116;
			7235: Pixel = 205;
			7236: Pixel = 182;
			7237: Pixel = 175;
			7238: Pixel = 153;
			7239: Pixel = 150;
			7240: Pixel = 137;
			7241: Pixel = 136;
			7242: Pixel = 120;
			7243: Pixel = 111;
			7244: Pixel = 105;
			7245: Pixel = 102;
			7246: Pixel = 129;
			7247: Pixel = 144;
			7248: Pixel = 135;
			7249: Pixel = 133;
			7250: Pixel = 133;
			7251: Pixel = 117;
			7252: Pixel = 122;
			7253: Pixel = 144;
			7254: Pixel = 145;
			7255: Pixel = 145;
			7256: Pixel = 137;
			7257: Pixel = 140;
			7258: Pixel = 132;
			7259: Pixel = 141;
			7260: Pixel = 152;
			7261: Pixel = 143;
			7262: Pixel = 140;
			7263: Pixel = 159;
			7264: Pixel = 158;
			7265: Pixel = 154;
			7266: Pixel = 158;
			7267: Pixel = 156;
			7268: Pixel = 158;
			7269: Pixel = 155;
			7270: Pixel = 153;
			7271: Pixel = 163;
			7272: Pixel = 171;
			7273: Pixel = 167;
			7274: Pixel = 152;
			7275: Pixel = 150;
			7276: Pixel = 160;
			7277: Pixel = 168;
			7278: Pixel = 163;
			7279: Pixel = 167;
			7280: Pixel = 162;
			7281: Pixel = 167;
			7282: Pixel = 168;
			7283: Pixel = 165;
			7284: Pixel = 163;
			7285: Pixel = 160;
			7286: Pixel = 165;
			7287: Pixel = 167;
			7288: Pixel = 163;
			7289: Pixel = 157;
			7290: Pixel = 152;
			7291: Pixel = 173;
			7292: Pixel = 189;
			7293: Pixel = 180;
			7294: Pixel = 179;
			7295: Pixel = 192;
			7296: Pixel = 200;
			7297: Pixel = 200;
			7298: Pixel = 193;
			7299: Pixel = 190;
			7300: Pixel = 191;
			7301: Pixel = 192;
			7302: Pixel = 195;
			7303: Pixel = 194;
			7304: Pixel = 197;
			7305: Pixel = 201;
			7306: Pixel = 202;
			7307: Pixel = 202;
			7308: Pixel = 201;
			7309: Pixel = 203;
			7310: Pixel = 206;
			7311: Pixel = 211;
			7312: Pixel = 196;
			7313: Pixel = 152;
			7314: Pixel = 169;
			7315: Pixel = 156;
			7316: Pixel = 159;
			7317: Pixel = 158;
			7318: Pixel = 176;
			7319: Pixel = 202;
			7320: Pixel = 55;
			7321: Pixel = 40;
			7322: Pixel = 48;
			7323: Pixel = 48;
			7324: Pixel = 49;
			7325: Pixel = 48;
			7326: Pixel = 49;
			7327: Pixel = 51;
			7328: Pixel = 49;
			7329: Pixel = 66;
			7330: Pixel = 117;
			7331: Pixel = 155;
			7332: Pixel = 147;
			7333: Pixel = 144;
			7334: Pixel = 154;
			7335: Pixel = 159;
			7336: Pixel = 160;
			7337: Pixel = 159;
			7338: Pixel = 157;
			7339: Pixel = 156;
			7340: Pixel = 156;
			7341: Pixel = 157;
			7342: Pixel = 157;
			7343: Pixel = 157;
			7344: Pixel = 156;
			7345: Pixel = 157;
			7346: Pixel = 156;
			7347: Pixel = 156;
			7348: Pixel = 156;
			7349: Pixel = 156;
			7350: Pixel = 95;
			7351: Pixel = 97;
			7352: Pixel = 97;
			7353: Pixel = 95;
			7354: Pixel = 96;
			7355: Pixel = 96;
			7356: Pixel = 100;
			7357: Pixel = 112;
			7358: Pixel = 132;
			7359: Pixel = 149;
			7360: Pixel = 162;
			7361: Pixel = 170;
			7362: Pixel = 171;
			7363: Pixel = 172;
			7364: Pixel = 172;
			7365: Pixel = 168;
			7366: Pixel = 157;
			7367: Pixel = 138;
			7368: Pixel = 106;
			7369: Pixel = 77;
			7370: Pixel = 77;
			7371: Pixel = 87;
			7372: Pixel = 94;
			7373: Pixel = 96;
			7374: Pixel = 98;
			7375: Pixel = 96;
			7376: Pixel = 96;
			7377: Pixel = 97;
			7378: Pixel = 98;
			7379: Pixel = 98;
			7380: Pixel = 97;
			7381: Pixel = 99;
			7382: Pixel = 99;
			7383: Pixel = 79;
			7384: Pixel = 124;
			7385: Pixel = 212;
			7386: Pixel = 190;
			7387: Pixel = 181;
			7388: Pixel = 167;
			7389: Pixel = 158;
			7390: Pixel = 144;
			7391: Pixel = 144;
			7392: Pixel = 131;
			7393: Pixel = 109;
			7394: Pixel = 94;
			7395: Pixel = 127;
			7396: Pixel = 137;
			7397: Pixel = 128;
			7398: Pixel = 133;
			7399: Pixel = 136;
			7400: Pixel = 119;
			7401: Pixel = 121;
			7402: Pixel = 140;
			7403: Pixel = 141;
			7404: Pixel = 144;
			7405: Pixel = 141;
			7406: Pixel = 136;
			7407: Pixel = 123;
			7408: Pixel = 137;
			7409: Pixel = 154;
			7410: Pixel = 140;
			7411: Pixel = 137;
			7412: Pixel = 159;
			7413: Pixel = 161;
			7414: Pixel = 157;
			7415: Pixel = 146;
			7416: Pixel = 152;
			7417: Pixel = 159;
			7418: Pixel = 157;
			7419: Pixel = 144;
			7420: Pixel = 134;
			7421: Pixel = 135;
			7422: Pixel = 118;
			7423: Pixel = 147;
			7424: Pixel = 162;
			7425: Pixel = 165;
			7426: Pixel = 161;
			7427: Pixel = 160;
			7428: Pixel = 162;
			7429: Pixel = 163;
			7430: Pixel = 167;
			7431: Pixel = 159;
			7432: Pixel = 161;
			7433: Pixel = 168;
			7434: Pixel = 166;
			7435: Pixel = 160;
			7436: Pixel = 161;
			7437: Pixel = 155;
			7438: Pixel = 149;
			7439: Pixel = 163;
			7440: Pixel = 185;
			7441: Pixel = 181;
			7442: Pixel = 178;
			7443: Pixel = 184;
			7444: Pixel = 201;
			7445: Pixel = 199;
			7446: Pixel = 189;
			7447: Pixel = 185;
			7448: Pixel = 183;
			7449: Pixel = 188;
			7450: Pixel = 193;
			7451: Pixel = 194;
			7452: Pixel = 196;
			7453: Pixel = 198;
			7454: Pixel = 201;
			7455: Pixel = 203;
			7456: Pixel = 203;
			7457: Pixel = 202;
			7458: Pixel = 202;
			7459: Pixel = 205;
			7460: Pixel = 209;
			7461: Pixel = 212;
			7462: Pixel = 164;
			7463: Pixel = 162;
			7464: Pixel = 157;
			7465: Pixel = 146;
			7466: Pixel = 126;
			7467: Pixel = 129;
			7468: Pixel = 211;
			7469: Pixel = 154;
			7470: Pixel = 28;
			7471: Pixel = 46;
			7472: Pixel = 53;
			7473: Pixel = 52;
			7474: Pixel = 50;
			7475: Pixel = 54;
			7476: Pixel = 61;
			7477: Pixel = 51;
			7478: Pixel = 51;
			7479: Pixel = 84;
			7480: Pixel = 144;
			7481: Pixel = 152;
			7482: Pixel = 144;
			7483: Pixel = 149;
			7484: Pixel = 158;
			7485: Pixel = 159;
			7486: Pixel = 158;
			7487: Pixel = 157;
			7488: Pixel = 156;
			7489: Pixel = 155;
			7490: Pixel = 156;
			7491: Pixel = 157;
			7492: Pixel = 157;
			7493: Pixel = 156;
			7494: Pixel = 156;
			7495: Pixel = 156;
			7496: Pixel = 156;
			7497: Pixel = 156;
			7498: Pixel = 156;
			7499: Pixel = 155;
			7500: Pixel = 97;
			7501: Pixel = 98;
			7502: Pixel = 97;
			7503: Pixel = 97;
			7504: Pixel = 97;
			7505: Pixel = 100;
			7506: Pixel = 105;
			7507: Pixel = 111;
			7508: Pixel = 131;
			7509: Pixel = 149;
			7510: Pixel = 162;
			7511: Pixel = 170;
			7512: Pixel = 172;
			7513: Pixel = 172;
			7514: Pixel = 171;
			7515: Pixel = 169;
			7516: Pixel = 158;
			7517: Pixel = 138;
			7518: Pixel = 102;
			7519: Pixel = 77;
			7520: Pixel = 75;
			7521: Pixel = 86;
			7522: Pixel = 94;
			7523: Pixel = 97;
			7524: Pixel = 98;
			7525: Pixel = 95;
			7526: Pixel = 94;
			7527: Pixel = 97;
			7528: Pixel = 97;
			7529: Pixel = 97;
			7530: Pixel = 99;
			7531: Pixel = 99;
			7532: Pixel = 97;
			7533: Pixel = 77;
			7534: Pixel = 122;
			7535: Pixel = 216;
			7536: Pixel = 194;
			7537: Pixel = 183;
			7538: Pixel = 167;
			7539: Pixel = 161;
			7540: Pixel = 152;
			7541: Pixel = 152;
			7542: Pixel = 145;
			7543: Pixel = 108;
			7544: Pixel = 109;
			7545: Pixel = 132;
			7546: Pixel = 131;
			7547: Pixel = 128;
			7548: Pixel = 136;
			7549: Pixel = 115;
			7550: Pixel = 121;
			7551: Pixel = 140;
			7552: Pixel = 143;
			7553: Pixel = 137;
			7554: Pixel = 141;
			7555: Pixel = 128;
			7556: Pixel = 125;
			7557: Pixel = 137;
			7558: Pixel = 143;
			7559: Pixel = 141;
			7560: Pixel = 135;
			7561: Pixel = 147;
			7562: Pixel = 155;
			7563: Pixel = 137;
			7564: Pixel = 117;
			7565: Pixel = 121;
			7566: Pixel = 111;
			7567: Pixel = 108;
			7568: Pixel = 129;
			7569: Pixel = 133;
			7570: Pixel = 133;
			7571: Pixel = 151;
			7572: Pixel = 110;
			7573: Pixel = 118;
			7574: Pixel = 153;
			7575: Pixel = 155;
			7576: Pixel = 164;
			7577: Pixel = 156;
			7578: Pixel = 152;
			7579: Pixel = 152;
			7580: Pixel = 161;
			7581: Pixel = 165;
			7582: Pixel = 156;
			7583: Pixel = 127;
			7584: Pixel = 136;
			7585: Pixel = 163;
			7586: Pixel = 148;
			7587: Pixel = 144;
			7588: Pixel = 173;
			7589: Pixel = 188;
			7590: Pixel = 175;
			7591: Pixel = 181;
			7592: Pixel = 195;
			7593: Pixel = 199;
			7594: Pixel = 197;
			7595: Pixel = 190;
			7596: Pixel = 188;
			7597: Pixel = 191;
			7598: Pixel = 191;
			7599: Pixel = 194;
			7600: Pixel = 197;
			7601: Pixel = 198;
			7602: Pixel = 198;
			7603: Pixel = 200;
			7604: Pixel = 202;
			7605: Pixel = 203;
			7606: Pixel = 203;
			7607: Pixel = 203;
			7608: Pixel = 203;
			7609: Pixel = 206;
			7610: Pixel = 215;
			7611: Pixel = 191;
			7612: Pixel = 161;
			7613: Pixel = 146;
			7614: Pixel = 107;
			7615: Pixel = 90;
			7616: Pixel = 102;
			7617: Pixel = 170;
			7618: Pixel = 228;
			7619: Pixel = 88;
			7620: Pixel = 25;
			7621: Pixel = 45;
			7622: Pixel = 50;
			7623: Pixel = 48;
			7624: Pixel = 46;
			7625: Pixel = 52;
			7626: Pixel = 55;
			7627: Pixel = 52;
			7628: Pixel = 59;
			7629: Pixel = 115;
			7630: Pixel = 155;
			7631: Pixel = 147;
			7632: Pixel = 146;
			7633: Pixel = 155;
			7634: Pixel = 159;
			7635: Pixel = 160;
			7636: Pixel = 158;
			7637: Pixel = 157;
			7638: Pixel = 156;
			7639: Pixel = 155;
			7640: Pixel = 155;
			7641: Pixel = 156;
			7642: Pixel = 155;
			7643: Pixel = 155;
			7644: Pixel = 155;
			7645: Pixel = 155;
			7646: Pixel = 156;
			7647: Pixel = 155;
			7648: Pixel = 154;
			7649: Pixel = 154;
			7650: Pixel = 98;
			7651: Pixel = 98;
			7652: Pixel = 97;
			7653: Pixel = 97;
			7654: Pixel = 99;
			7655: Pixel = 99;
			7656: Pixel = 103;
			7657: Pixel = 112;
			7658: Pixel = 133;
			7659: Pixel = 149;
			7660: Pixel = 162;
			7661: Pixel = 170;
			7662: Pixel = 172;
			7663: Pixel = 173;
			7664: Pixel = 172;
			7665: Pixel = 170;
			7666: Pixel = 160;
			7667: Pixel = 137;
			7668: Pixel = 104;
			7669: Pixel = 75;
			7670: Pixel = 75;
			7671: Pixel = 86;
			7672: Pixel = 92;
			7673: Pixel = 98;
			7674: Pixel = 97;
			7675: Pixel = 98;
			7676: Pixel = 99;
			7677: Pixel = 98;
			7678: Pixel = 99;
			7679: Pixel = 98;
			7680: Pixel = 99;
			7681: Pixel = 97;
			7682: Pixel = 96;
			7683: Pixel = 77;
			7684: Pixel = 119;
			7685: Pixel = 216;
			7686: Pixel = 196;
			7687: Pixel = 189;
			7688: Pixel = 170;
			7689: Pixel = 160;
			7690: Pixel = 150;
			7691: Pixel = 153;
			7692: Pixel = 148;
			7693: Pixel = 122;
			7694: Pixel = 120;
			7695: Pixel = 119;
			7696: Pixel = 123;
			7697: Pixel = 134;
			7698: Pixel = 116;
			7699: Pixel = 116;
			7700: Pixel = 138;
			7701: Pixel = 140;
			7702: Pixel = 137;
			7703: Pixel = 136;
			7704: Pixel = 125;
			7705: Pixel = 124;
			7706: Pixel = 131;
			7707: Pixel = 142;
			7708: Pixel = 137;
			7709: Pixel = 130;
			7710: Pixel = 149;
			7711: Pixel = 155;
			7712: Pixel = 133;
			7713: Pixel = 107;
			7714: Pixel = 137;
			7715: Pixel = 134;
			7716: Pixel = 118;
			7717: Pixel = 104;
			7718: Pixel = 90;
			7719: Pixel = 78;
			7720: Pixel = 143;
			7721: Pixel = 174;
			7722: Pixel = 159;
			7723: Pixel = 122;
			7724: Pixel = 119;
			7725: Pixel = 124;
			7726: Pixel = 116;
			7727: Pixel = 132;
			7728: Pixel = 148;
			7729: Pixel = 134;
			7730: Pixel = 118;
			7731: Pixel = 117;
			7732: Pixel = 109;
			7733: Pixel = 102;
			7734: Pixel = 61;
			7735: Pixel = 124;
			7736: Pixel = 155;
			7737: Pixel = 178;
			7738: Pixel = 175;
			7739: Pixel = 164;
			7740: Pixel = 182;
			7741: Pixel = 200;
			7742: Pixel = 202;
			7743: Pixel = 193;
			7744: Pixel = 194;
			7745: Pixel = 194;
			7746: Pixel = 194;
			7747: Pixel = 191;
			7748: Pixel = 194;
			7749: Pixel = 196;
			7750: Pixel = 200;
			7751: Pixel = 200;
			7752: Pixel = 201;
			7753: Pixel = 201;
			7754: Pixel = 204;
			7755: Pixel = 203;
			7756: Pixel = 201;
			7757: Pixel = 201;
			7758: Pixel = 207;
			7759: Pixel = 217;
			7760: Pixel = 202;
			7761: Pixel = 159;
			7762: Pixel = 120;
			7763: Pixel = 86;
			7764: Pixel = 84;
			7765: Pixel = 99;
			7766: Pixel = 150;
			7767: Pixel = 221;
			7768: Pixel = 172;
			7769: Pixel = 34;
			7770: Pixel = 41;
			7771: Pixel = 46;
			7772: Pixel = 49;
			7773: Pixel = 45;
			7774: Pixel = 44;
			7775: Pixel = 54;
			7776: Pixel = 54;
			7777: Pixel = 49;
			7778: Pixel = 81;
			7779: Pixel = 141;
			7780: Pixel = 151;
			7781: Pixel = 145;
			7782: Pixel = 151;
			7783: Pixel = 161;
			7784: Pixel = 159;
			7785: Pixel = 158;
			7786: Pixel = 159;
			7787: Pixel = 157;
			7788: Pixel = 156;
			7789: Pixel = 156;
			7790: Pixel = 156;
			7791: Pixel = 156;
			7792: Pixel = 155;
			7793: Pixel = 154;
			7794: Pixel = 154;
			7795: Pixel = 155;
			7796: Pixel = 154;
			7797: Pixel = 154;
			7798: Pixel = 152;
			7799: Pixel = 153;
			7800: Pixel = 99;
			7801: Pixel = 99;
			7802: Pixel = 99;
			7803: Pixel = 98;
			7804: Pixel = 100;
			7805: Pixel = 102;
			7806: Pixel = 105;
			7807: Pixel = 117;
			7808: Pixel = 135;
			7809: Pixel = 151;
			7810: Pixel = 163;
			7811: Pixel = 172;
			7812: Pixel = 172;
			7813: Pixel = 174;
			7814: Pixel = 173;
			7815: Pixel = 171;
			7816: Pixel = 159;
			7817: Pixel = 138;
			7818: Pixel = 104;
			7819: Pixel = 75;
			7820: Pixel = 74;
			7821: Pixel = 84;
			7822: Pixel = 93;
			7823: Pixel = 95;
			7824: Pixel = 96;
			7825: Pixel = 101;
			7826: Pixel = 99;
			7827: Pixel = 100;
			7828: Pixel = 99;
			7829: Pixel = 98;
			7830: Pixel = 99;
			7831: Pixel = 99;
			7832: Pixel = 96;
			7833: Pixel = 80;
			7834: Pixel = 113;
			7835: Pixel = 215;
			7836: Pixel = 197;
			7837: Pixel = 193;
			7838: Pixel = 185;
			7839: Pixel = 161;
			7840: Pixel = 135;
			7841: Pixel = 143;
			7842: Pixel = 152;
			7843: Pixel = 114;
			7844: Pixel = 111;
			7845: Pixel = 121;
			7846: Pixel = 124;
			7847: Pixel = 110;
			7848: Pixel = 113;
			7849: Pixel = 135;
			7850: Pixel = 139;
			7851: Pixel = 136;
			7852: Pixel = 137;
			7853: Pixel = 123;
			7854: Pixel = 123;
			7855: Pixel = 131;
			7856: Pixel = 136;
			7857: Pixel = 128;
			7858: Pixel = 131;
			7859: Pixel = 143;
			7860: Pixel = 143;
			7861: Pixel = 134;
			7862: Pixel = 122;
			7863: Pixel = 149;
			7864: Pixel = 124;
			7865: Pixel = 102;
			7866: Pixel = 100;
			7867: Pixel = 86;
			7868: Pixel = 80;
			7869: Pixel = 73;
			7870: Pixel = 135;
			7871: Pixel = 158;
			7872: Pixel = 145;
			7873: Pixel = 126;
			7874: Pixel = 106;
			7875: Pixel = 92;
			7876: Pixel = 80;
			7877: Pixel = 94;
			7878: Pixel = 77;
			7879: Pixel = 77;
			7880: Pixel = 66;
			7881: Pixel = 51;
			7882: Pixel = 45;
			7883: Pixel = 51;
			7884: Pixel = 30;
			7885: Pixel = 109;
			7886: Pixel = 190;
			7887: Pixel = 159;
			7888: Pixel = 166;
			7889: Pixel = 191;
			7890: Pixel = 199;
			7891: Pixel = 195;
			7892: Pixel = 194;
			7893: Pixel = 192;
			7894: Pixel = 196;
			7895: Pixel = 195;
			7896: Pixel = 192;
			7897: Pixel = 192;
			7898: Pixel = 195;
			7899: Pixel = 198;
			7900: Pixel = 200;
			7901: Pixel = 200;
			7902: Pixel = 200;
			7903: Pixel = 200;
			7904: Pixel = 204;
			7905: Pixel = 202;
			7906: Pixel = 209;
			7907: Pixel = 212;
			7908: Pixel = 199;
			7909: Pixel = 165;
			7910: Pixel = 125;
			7911: Pixel = 94;
			7912: Pixel = 80;
			7913: Pixel = 87;
			7914: Pixel = 98;
			7915: Pixel = 139;
			7916: Pixel = 199;
			7917: Pixel = 216;
			7918: Pixel = 73;
			7919: Pixel = 32;
			7920: Pixel = 49;
			7921: Pixel = 50;
			7922: Pixel = 47;
			7923: Pixel = 44;
			7924: Pixel = 47;
			7925: Pixel = 54;
			7926: Pixel = 45;
			7927: Pixel = 52;
			7928: Pixel = 116;
			7929: Pixel = 152;
			7930: Pixel = 145;
			7931: Pixel = 144;
			7932: Pixel = 158;
			7933: Pixel = 160;
			7934: Pixel = 160;
			7935: Pixel = 159;
			7936: Pixel = 158;
			7937: Pixel = 159;
			7938: Pixel = 157;
			7939: Pixel = 155;
			7940: Pixel = 156;
			7941: Pixel = 155;
			7942: Pixel = 154;
			7943: Pixel = 155;
			7944: Pixel = 154;
			7945: Pixel = 154;
			7946: Pixel = 153;
			7947: Pixel = 154;
			7948: Pixel = 154;
			7949: Pixel = 153;
			7950: Pixel = 98;
			7951: Pixel = 102;
			7952: Pixel = 102;
			7953: Pixel = 98;
			7954: Pixel = 98;
			7955: Pixel = 102;
			7956: Pixel = 108;
			7957: Pixel = 115;
			7958: Pixel = 134;
			7959: Pixel = 152;
			7960: Pixel = 165;
			7961: Pixel = 171;
			7962: Pixel = 172;
			7963: Pixel = 172;
			7964: Pixel = 173;
			7965: Pixel = 171;
			7966: Pixel = 159;
			7967: Pixel = 140;
			7968: Pixel = 104;
			7969: Pixel = 74;
			7970: Pixel = 76;
			7971: Pixel = 85;
			7972: Pixel = 94;
			7973: Pixel = 96;
			7974: Pixel = 98;
			7975: Pixel = 97;
			7976: Pixel = 98;
			7977: Pixel = 100;
			7978: Pixel = 98;
			7979: Pixel = 99;
			7980: Pixel = 99;
			7981: Pixel = 100;
			7982: Pixel = 98;
			7983: Pixel = 87;
			7984: Pixel = 94;
			7985: Pixel = 203;
			7986: Pixel = 202;
			7987: Pixel = 199;
			7988: Pixel = 192;
			7989: Pixel = 160;
			7990: Pixel = 123;
			7991: Pixel = 126;
			7992: Pixel = 129;
			7993: Pixel = 110;
			7994: Pixel = 111;
			7995: Pixel = 123;
			7996: Pixel = 113;
			7997: Pixel = 106;
			7998: Pixel = 130;
			7999: Pixel = 138;
			8000: Pixel = 133;
			8001: Pixel = 135;
			8002: Pixel = 121;
			8003: Pixel = 127;
			8004: Pixel = 134;
			8005: Pixel = 132;
			8006: Pixel = 132;
			8007: Pixel = 126;
			8008: Pixel = 140;
			8009: Pixel = 144;
			8010: Pixel = 131;
			8011: Pixel = 110;
			8012: Pixel = 137;
			8013: Pixel = 128;
			8014: Pixel = 108;
			8015: Pixel = 120;
			8016: Pixel = 109;
			8017: Pixel = 127;
			8018: Pixel = 102;
			8019: Pixel = 86;
			8020: Pixel = 98;
			8021: Pixel = 111;
			8022: Pixel = 115;
			8023: Pixel = 84;
			8024: Pixel = 60;
			8025: Pixel = 69;
			8026: Pixel = 96;
			8027: Pixel = 81;
			8028: Pixel = 67;
			8029: Pixel = 66;
			8030: Pixel = 42;
			8031: Pixel = 40;
			8032: Pixel = 40;
			8033: Pixel = 47;
			8034: Pixel = 125;
			8035: Pixel = 168;
			8036: Pixel = 148;
			8037: Pixel = 180;
			8038: Pixel = 205;
			8039: Pixel = 200;
			8040: Pixel = 195;
			8041: Pixel = 194;
			8042: Pixel = 192;
			8043: Pixel = 194;
			8044: Pixel = 195;
			8045: Pixel = 194;
			8046: Pixel = 191;
			8047: Pixel = 194;
			8048: Pixel = 195;
			8049: Pixel = 197;
			8050: Pixel = 198;
			8051: Pixel = 200;
			8052: Pixel = 197;
			8053: Pixel = 200;
			8054: Pixel = 208;
			8055: Pixel = 211;
			8056: Pixel = 187;
			8057: Pixel = 141;
			8058: Pixel = 104;
			8059: Pixel = 85;
			8060: Pixel = 88;
			8061: Pixel = 87;
			8062: Pixel = 90;
			8063: Pixel = 108;
			8064: Pixel = 143;
			8065: Pixel = 192;
			8066: Pixel = 207;
			8067: Pixel = 115;
			8068: Pixel = 37;
			8069: Pixel = 46;
			8070: Pixel = 51;
			8071: Pixel = 50;
			8072: Pixel = 50;
			8073: Pixel = 47;
			8074: Pixel = 53;
			8075: Pixel = 51;
			8076: Pixel = 37;
			8077: Pixel = 69;
			8078: Pixel = 141;
			8079: Pixel = 149;
			8080: Pixel = 142;
			8081: Pixel = 152;
			8082: Pixel = 163;
			8083: Pixel = 160;
			8084: Pixel = 160;
			8085: Pixel = 160;
			8086: Pixel = 159;
			8087: Pixel = 159;
			8088: Pixel = 157;
			8089: Pixel = 157;
			8090: Pixel = 156;
			8091: Pixel = 154;
			8092: Pixel = 153;
			8093: Pixel = 154;
			8094: Pixel = 155;
			8095: Pixel = 154;
			8096: Pixel = 154;
			8097: Pixel = 153;
			8098: Pixel = 153;
			8099: Pixel = 153;
			8100: Pixel = 100;
			8101: Pixel = 102;
			8102: Pixel = 103;
			8103: Pixel = 99;
			8104: Pixel = 95;
			8105: Pixel = 104;
			8106: Pixel = 107;
			8107: Pixel = 116;
			8108: Pixel = 134;
			8109: Pixel = 151;
			8110: Pixel = 165;
			8111: Pixel = 172;
			8112: Pixel = 170;
			8113: Pixel = 172;
			8114: Pixel = 173;
			8115: Pixel = 170;
			8116: Pixel = 160;
			8117: Pixel = 139;
			8118: Pixel = 103;
			8119: Pixel = 75;
			8120: Pixel = 77;
			8121: Pixel = 86;
			8122: Pixel = 94;
			8123: Pixel = 95;
			8124: Pixel = 98;
			8125: Pixel = 98;
			8126: Pixel = 98;
			8127: Pixel = 101;
			8128: Pixel = 99;
			8129: Pixel = 99;
			8130: Pixel = 99;
			8131: Pixel = 97;
			8132: Pixel = 95;
			8133: Pixel = 90;
			8134: Pixel = 79;
			8135: Pixel = 186;
			8136: Pixel = 211;
			8137: Pixel = 199;
			8138: Pixel = 196;
			8139: Pixel = 162;
			8140: Pixel = 117;
			8141: Pixel = 128;
			8142: Pixel = 143;
			8143: Pixel = 126;
			8144: Pixel = 122;
			8145: Pixel = 109;
			8146: Pixel = 108;
			8147: Pixel = 126;
			8148: Pixel = 138;
			8149: Pixel = 137;
			8150: Pixel = 133;
			8151: Pixel = 121;
			8152: Pixel = 121;
			8153: Pixel = 130;
			8154: Pixel = 136;
			8155: Pixel = 131;
			8156: Pixel = 123;
			8157: Pixel = 137;
			8158: Pixel = 140;
			8159: Pixel = 130;
			8160: Pixel = 114;
			8161: Pixel = 131;
			8162: Pixel = 132;
			8163: Pixel = 112;
			8164: Pixel = 126;
			8165: Pixel = 113;
			8166: Pixel = 93;
			8167: Pixel = 79;
			8168: Pixel = 63;
			8169: Pixel = 59;
			8170: Pixel = 69;
			8171: Pixel = 102;
			8172: Pixel = 111;
			8173: Pixel = 94;
			8174: Pixel = 99;
			8175: Pixel = 106;
			8176: Pixel = 87;
			8177: Pixel = 59;
			8178: Pixel = 73;
			8179: Pixel = 74;
			8180: Pixel = 42;
			8181: Pixel = 32;
			8182: Pixel = 41;
			8183: Pixel = 142;
			8184: Pixel = 162;
			8185: Pixel = 141;
			8186: Pixel = 184;
			8187: Pixel = 194;
			8188: Pixel = 194;
			8189: Pixel = 195;
			8190: Pixel = 194;
			8191: Pixel = 192;
			8192: Pixel = 192;
			8193: Pixel = 190;
			8194: Pixel = 193;
			8195: Pixel = 193;
			8196: Pixel = 191;
			8197: Pixel = 192;
			8198: Pixel = 194;
			8199: Pixel = 196;
			8200: Pixel = 197;
			8201: Pixel = 200;
			8202: Pixel = 202;
			8203: Pixel = 213;
			8204: Pixel = 202;
			8205: Pixel = 139;
			8206: Pixel = 91;
			8207: Pixel = 84;
			8208: Pixel = 83;
			8209: Pixel = 85;
			8210: Pixel = 96;
			8211: Pixel = 106;
			8212: Pixel = 127;
			8213: Pixel = 164;
			8214: Pixel = 200;
			8215: Pixel = 188;
			8216: Pixel = 72;
			8217: Pixel = 35;
			8218: Pixel = 43;
			8219: Pixel = 50;
			8220: Pixel = 50;
			8221: Pixel = 47;
			8222: Pixel = 47;
			8223: Pixel = 50;
			8224: Pixel = 56;
			8225: Pixel = 49;
			8226: Pixel = 42;
			8227: Pixel = 102;
			8228: Pixel = 151;
			8229: Pixel = 145;
			8230: Pixel = 145;
			8231: Pixel = 160;
			8232: Pixel = 164;
			8233: Pixel = 162;
			8234: Pixel = 160;
			8235: Pixel = 160;
			8236: Pixel = 160;
			8237: Pixel = 159;
			8238: Pixel = 158;
			8239: Pixel = 157;
			8240: Pixel = 155;
			8241: Pixel = 156;
			8242: Pixel = 156;
			8243: Pixel = 154;
			8244: Pixel = 153;
			8245: Pixel = 154;
			8246: Pixel = 154;
			8247: Pixel = 153;
			8248: Pixel = 153;
			8249: Pixel = 152;
			8250: Pixel = 105;
			8251: Pixel = 104;
			8252: Pixel = 102;
			8253: Pixel = 98;
			8254: Pixel = 98;
			8255: Pixel = 101;
			8256: Pixel = 106;
			8257: Pixel = 114;
			8258: Pixel = 135;
			8259: Pixel = 149;
			8260: Pixel = 163;
			8261: Pixel = 171;
			8262: Pixel = 171;
			8263: Pixel = 171;
			8264: Pixel = 172;
			8265: Pixel = 169;
			8266: Pixel = 160;
			8267: Pixel = 139;
			8268: Pixel = 104;
			8269: Pixel = 77;
			8270: Pixel = 76;
			8271: Pixel = 85;
			8272: Pixel = 93;
			8273: Pixel = 95;
			8274: Pixel = 97;
			8275: Pixel = 97;
			8276: Pixel = 97;
			8277: Pixel = 101;
			8278: Pixel = 98;
			8279: Pixel = 97;
			8280: Pixel = 100;
			8281: Pixel = 96;
			8282: Pixel = 96;
			8283: Pixel = 97;
			8284: Pixel = 74;
			8285: Pixel = 158;
			8286: Pixel = 213;
			8287: Pixel = 197;
			8288: Pixel = 198;
			8289: Pixel = 160;
			8290: Pixel = 129;
			8291: Pixel = 142;
			8292: Pixel = 147;
			8293: Pixel = 139;
			8294: Pixel = 115;
			8295: Pixel = 102;
			8296: Pixel = 119;
			8297: Pixel = 134;
			8298: Pixel = 135;
			8299: Pixel = 135;
			8300: Pixel = 120;
			8301: Pixel = 123;
			8302: Pixel = 127;
			8303: Pixel = 134;
			8304: Pixel = 130;
			8305: Pixel = 123;
			8306: Pixel = 138;
			8307: Pixel = 137;
			8308: Pixel = 133;
			8309: Pixel = 107;
			8310: Pixel = 127;
			8311: Pixel = 138;
			8312: Pixel = 119;
			8313: Pixel = 91;
			8314: Pixel = 81;
			8315: Pixel = 85;
			8316: Pixel = 74;
			8317: Pixel = 54;
			8318: Pixel = 53;
			8319: Pixel = 58;
			8320: Pixel = 99;
			8321: Pixel = 116;
			8322: Pixel = 92;
			8323: Pixel = 61;
			8324: Pixel = 91;
			8325: Pixel = 98;
			8326: Pixel = 92;
			8327: Pixel = 68;
			8328: Pixel = 65;
			8329: Pixel = 73;
			8330: Pixel = 17;
			8331: Pixel = 60;
			8332: Pixel = 159;
			8333: Pixel = 150;
			8334: Pixel = 127;
			8335: Pixel = 186;
			8336: Pixel = 195;
			8337: Pixel = 179;
			8338: Pixel = 183;
			8339: Pixel = 192;
			8340: Pixel = 191;
			8341: Pixel = 191;
			8342: Pixel = 188;
			8343: Pixel = 187;
			8344: Pixel = 191;
			8345: Pixel = 190;
			8346: Pixel = 190;
			8347: Pixel = 192;
			8348: Pixel = 194;
			8349: Pixel = 194;
			8350: Pixel = 198;
			8351: Pixel = 206;
			8352: Pixel = 196;
			8353: Pixel = 152;
			8354: Pixel = 134;
			8355: Pixel = 103;
			8356: Pixel = 90;
			8357: Pixel = 90;
			8358: Pixel = 94;
			8359: Pixel = 110;
			8360: Pixel = 137;
			8361: Pixel = 158;
			8362: Pixel = 168;
			8363: Pixel = 191;
			8364: Pixel = 200;
			8365: Pixel = 82;
			8366: Pixel = 33;
			8367: Pixel = 49;
			8368: Pixel = 49;
			8369: Pixel = 54;
			8370: Pixel = 50;
			8371: Pixel = 44;
			8372: Pixel = 44;
			8373: Pixel = 53;
			8374: Pixel = 61;
			8375: Pixel = 53;
			8376: Pixel = 66;
			8377: Pixel = 133;
			8378: Pixel = 151;
			8379: Pixel = 143;
			8380: Pixel = 153;
			8381: Pixel = 165;
			8382: Pixel = 163;
			8383: Pixel = 161;
			8384: Pixel = 161;
			8385: Pixel = 160;
			8386: Pixel = 160;
			8387: Pixel = 159;
			8388: Pixel = 159;
			8389: Pixel = 157;
			8390: Pixel = 158;
			8391: Pixel = 156;
			8392: Pixel = 155;
			8393: Pixel = 156;
			8394: Pixel = 155;
			8395: Pixel = 154;
			8396: Pixel = 154;
			8397: Pixel = 154;
			8398: Pixel = 153;
			8399: Pixel = 151;
			8400: Pixel = 106;
			8401: Pixel = 105;
			8402: Pixel = 103;
			8403: Pixel = 102;
			8404: Pixel = 101;
			8405: Pixel = 99;
			8406: Pixel = 103;
			8407: Pixel = 114;
			8408: Pixel = 134;
			8409: Pixel = 150;
			8410: Pixel = 162;
			8411: Pixel = 169;
			8412: Pixel = 170;
			8413: Pixel = 170;
			8414: Pixel = 170;
			8415: Pixel = 169;
			8416: Pixel = 159;
			8417: Pixel = 141;
			8418: Pixel = 105;
			8419: Pixel = 77;
			8420: Pixel = 75;
			8421: Pixel = 84;
			8422: Pixel = 91;
			8423: Pixel = 95;
			8424: Pixel = 96;
			8425: Pixel = 98;
			8426: Pixel = 97;
			8427: Pixel = 99;
			8428: Pixel = 98;
			8429: Pixel = 98;
			8430: Pixel = 99;
			8431: Pixel = 99;
			8432: Pixel = 100;
			8433: Pixel = 99;
			8434: Pixel = 77;
			8435: Pixel = 115;
			8436: Pixel = 213;
			8437: Pixel = 194;
			8438: Pixel = 194;
			8439: Pixel = 178;
			8440: Pixel = 140;
			8441: Pixel = 132;
			8442: Pixel = 146;
			8443: Pixel = 136;
			8444: Pixel = 102;
			8445: Pixel = 116;
			8446: Pixel = 133;
			8447: Pixel = 135;
			8448: Pixel = 134;
			8449: Pixel = 116;
			8450: Pixel = 120;
			8451: Pixel = 129;
			8452: Pixel = 126;
			8453: Pixel = 131;
			8454: Pixel = 121;
			8455: Pixel = 131;
			8456: Pixel = 141;
			8457: Pixel = 138;
			8458: Pixel = 135;
			8459: Pixel = 109;
			8460: Pixel = 135;
			8461: Pixel = 102;
			8462: Pixel = 67;
			8463: Pixel = 68;
			8464: Pixel = 88;
			8465: Pixel = 68;
			8466: Pixel = 57;
			8467: Pixel = 53;
			8468: Pixel = 45;
			8469: Pixel = 87;
			8470: Pixel = 128;
			8471: Pixel = 92;
			8472: Pixel = 41;
			8473: Pixel = 58;
			8474: Pixel = 95;
			8475: Pixel = 80;
			8476: Pixel = 86;
			8477: Pixel = 37;
			8478: Pixel = 68;
			8479: Pixel = 69;
			8480: Pixel = 63;
			8481: Pixel = 158;
			8482: Pixel = 142;
			8483: Pixel = 146;
			8484: Pixel = 195;
			8485: Pixel = 192;
			8486: Pixel = 180;
			8487: Pixel = 179;
			8488: Pixel = 186;
			8489: Pixel = 187;
			8490: Pixel = 187;
			8491: Pixel = 188;
			8492: Pixel = 185;
			8493: Pixel = 187;
			8494: Pixel = 189;
			8495: Pixel = 190;
			8496: Pixel = 191;
			8497: Pixel = 193;
			8498: Pixel = 193;
			8499: Pixel = 205;
			8500: Pixel = 200;
			8501: Pixel = 160;
			8502: Pixel = 100;
			8503: Pixel = 95;
			8504: Pixel = 127;
			8505: Pixel = 138;
			8506: Pixel = 123;
			8507: Pixel = 131;
			8508: Pixel = 152;
			8509: Pixel = 165;
			8510: Pixel = 169;
			8511: Pixel = 164;
			8512: Pixel = 183;
			8513: Pixel = 197;
			8514: Pixel = 81;
			8515: Pixel = 32;
			8516: Pixel = 49;
			8517: Pixel = 51;
			8518: Pixel = 55;
			8519: Pixel = 53;
			8520: Pixel = 50;
			8521: Pixel = 46;
			8522: Pixel = 43;
			8523: Pixel = 57;
			8524: Pixel = 55;
			8525: Pixel = 49;
			8526: Pixel = 97;
			8527: Pixel = 149;
			8528: Pixel = 146;
			8529: Pixel = 143;
			8530: Pixel = 161;
			8531: Pixel = 164;
			8532: Pixel = 164;
			8533: Pixel = 164;
			8534: Pixel = 163;
			8535: Pixel = 161;
			8536: Pixel = 162;
			8537: Pixel = 160;
			8538: Pixel = 159;
			8539: Pixel = 158;
			8540: Pixel = 158;
			8541: Pixel = 156;
			8542: Pixel = 154;
			8543: Pixel = 155;
			8544: Pixel = 154;
			8545: Pixel = 155;
			8546: Pixel = 155;
			8547: Pixel = 155;
			8548: Pixel = 152;
			8549: Pixel = 150;
			8550: Pixel = 108;
			8551: Pixel = 104;
			8552: Pixel = 103;
			8553: Pixel = 104;
			8554: Pixel = 99;
			8555: Pixel = 101;
			8556: Pixel = 103;
			8557: Pixel = 113;
			8558: Pixel = 132;
			8559: Pixel = 150;
			8560: Pixel = 162;
			8561: Pixel = 171;
			8562: Pixel = 170;
			8563: Pixel = 171;
			8564: Pixel = 171;
			8565: Pixel = 170;
			8566: Pixel = 159;
			8567: Pixel = 139;
			8568: Pixel = 107;
			8569: Pixel = 76;
			8570: Pixel = 76;
			8571: Pixel = 86;
			8572: Pixel = 92;
			8573: Pixel = 95;
			8574: Pixel = 95;
			8575: Pixel = 98;
			8576: Pixel = 99;
			8577: Pixel = 100;
			8578: Pixel = 99;
			8579: Pixel = 98;
			8580: Pixel = 97;
			8581: Pixel = 97;
			8582: Pixel = 100;
			8583: Pixel = 101;
			8584: Pixel = 87;
			8585: Pixel = 87;
			8586: Pixel = 201;
			8587: Pixel = 200;
			8588: Pixel = 195;
			8589: Pixel = 191;
			8590: Pixel = 165;
			8591: Pixel = 151;
			8592: Pixel = 150;
			8593: Pixel = 111;
			8594: Pixel = 112;
			8595: Pixel = 131;
			8596: Pixel = 138;
			8597: Pixel = 136;
			8598: Pixel = 109;
			8599: Pixel = 113;
			8600: Pixel = 128;
			8601: Pixel = 127;
			8602: Pixel = 128;
			8603: Pixel = 119;
			8604: Pixel = 122;
			8605: Pixel = 126;
			8606: Pixel = 112;
			8607: Pixel = 125;
			8608: Pixel = 146;
			8609: Pixel = 111;
			8610: Pixel = 90;
			8611: Pixel = 61;
			8612: Pixel = 71;
			8613: Pixel = 83;
			8614: Pixel = 54;
			8615: Pixel = 44;
			8616: Pixel = 55;
			8617: Pixel = 41;
			8618: Pixel = 58;
			8619: Pixel = 110;
			8620: Pixel = 86;
			8621: Pixel = 49;
			8622: Pixel = 61;
			8623: Pixel = 114;
			8624: Pixel = 96;
			8625: Pixel = 77;
			8626: Pixel = 47;
			8627: Pixel = 43;
			8628: Pixel = 70;
			8629: Pixel = 105;
			8630: Pixel = 160;
			8631: Pixel = 135;
			8632: Pixel = 150;
			8633: Pixel = 199;
			8634: Pixel = 192;
			8635: Pixel = 180;
			8636: Pixel = 179;
			8637: Pixel = 183;
			8638: Pixel = 184;
			8639: Pixel = 180;
			8640: Pixel = 180;
			8641: Pixel = 181;
			8642: Pixel = 183;
			8643: Pixel = 186;
			8644: Pixel = 190;
			8645: Pixel = 191;
			8646: Pixel = 191;
			8647: Pixel = 195;
			8648: Pixel = 205;
			8649: Pixel = 170;
			8650: Pixel = 97;
			8651: Pixel = 69;
			8652: Pixel = 106;
			8653: Pixel = 103;
			8654: Pixel = 117;
			8655: Pixel = 152;
			8656: Pixel = 167;
			8657: Pixel = 168;
			8658: Pixel = 169;
			8659: Pixel = 166;
			8660: Pixel = 168;
			8661: Pixel = 187;
			8662: Pixel = 204;
			8663: Pixel = 93;
			8664: Pixel = 28;
			8665: Pixel = 45;
			8666: Pixel = 49;
			8667: Pixel = 55;
			8668: Pixel = 54;
			8669: Pixel = 52;
			8670: Pixel = 48;
			8671: Pixel = 47;
			8672: Pixel = 50;
			8673: Pixel = 54;
			8674: Pixel = 44;
			8675: Pixel = 57;
			8676: Pixel = 127;
			8677: Pixel = 150;
			8678: Pixel = 142;
			8679: Pixel = 150;
			8680: Pixel = 165;
			8681: Pixel = 164;
			8682: Pixel = 164;
			8683: Pixel = 166;
			8684: Pixel = 163;
			8685: Pixel = 161;
			8686: Pixel = 162;
			8687: Pixel = 161;
			8688: Pixel = 158;
			8689: Pixel = 158;
			8690: Pixel = 158;
			8691: Pixel = 157;
			8692: Pixel = 156;
			8693: Pixel = 155;
			8694: Pixel = 155;
			8695: Pixel = 155;
			8696: Pixel = 154;
			8697: Pixel = 153;
			8698: Pixel = 153;
			8699: Pixel = 151;
			8700: Pixel = 105;
			8701: Pixel = 105;
			8702: Pixel = 104;
			8703: Pixel = 102;
			8704: Pixel = 100;
			8705: Pixel = 101;
			8706: Pixel = 101;
			8707: Pixel = 110;
			8708: Pixel = 131;
			8709: Pixel = 148;
			8710: Pixel = 163;
			8711: Pixel = 171;
			8712: Pixel = 171;
			8713: Pixel = 171;
			8714: Pixel = 171;
			8715: Pixel = 170;
			8716: Pixel = 159;
			8717: Pixel = 142;
			8718: Pixel = 109;
			8719: Pixel = 75;
			8720: Pixel = 74;
			8721: Pixel = 87;
			8722: Pixel = 91;
			8723: Pixel = 93;
			8724: Pixel = 96;
			8725: Pixel = 95;
			8726: Pixel = 97;
			8727: Pixel = 100;
			8728: Pixel = 96;
			8729: Pixel = 96;
			8730: Pixel = 98;
			8731: Pixel = 99;
			8732: Pixel = 104;
			8733: Pixel = 103;
			8734: Pixel = 98;
			8735: Pixel = 80;
			8736: Pixel = 159;
			8737: Pixel = 217;
			8738: Pixel = 201;
			8739: Pixel = 179;
			8740: Pixel = 168;
			8741: Pixel = 172;
			8742: Pixel = 133;
			8743: Pixel = 101;
			8744: Pixel = 127;
			8745: Pixel = 129;
			8746: Pixel = 135;
			8747: Pixel = 117;
			8748: Pixel = 116;
			8749: Pixel = 126;
			8750: Pixel = 126;
			8751: Pixel = 119;
			8752: Pixel = 122;
			8753: Pixel = 122;
			8754: Pixel = 140;
			8755: Pixel = 140;
			8756: Pixel = 110;
			8757: Pixel = 89;
			8758: Pixel = 98;
			8759: Pixel = 90;
			8760: Pixel = 61;
			8761: Pixel = 80;
			8762: Pixel = 81;
			8763: Pixel = 57;
			8764: Pixel = 53;
			8765: Pixel = 75;
			8766: Pixel = 44;
			8767: Pixel = 40;
			8768: Pixel = 88;
			8769: Pixel = 82;
			8770: Pixel = 46;
			8771: Pixel = 57;
			8772: Pixel = 95;
			8773: Pixel = 93;
			8774: Pixel = 103;
			8775: Pixel = 52;
			8776: Pixel = 94;
			8777: Pixel = 39;
			8778: Pixel = 122;
			8779: Pixel = 159;
			8780: Pixel = 121;
			8781: Pixel = 160;
			8782: Pixel = 199;
			8783: Pixel = 193;
			8784: Pixel = 187;
			8785: Pixel = 177;
			8786: Pixel = 180;
			8787: Pixel = 181;
			8788: Pixel = 181;
			8789: Pixel = 178;
			8790: Pixel = 177;
			8791: Pixel = 175;
			8792: Pixel = 180;
			8793: Pixel = 189;
			8794: Pixel = 191;
			8795: Pixel = 190;
			8796: Pixel = 193;
			8797: Pixel = 190;
			8798: Pixel = 136;
			8799: Pixel = 47;
			8800: Pixel = 84;
			8801: Pixel = 89;
			8802: Pixel = 128;
			8803: Pixel = 117;
			8804: Pixel = 115;
			8805: Pixel = 144;
			8806: Pixel = 159;
			8807: Pixel = 167;
			8808: Pixel = 169;
			8809: Pixel = 170;
			8810: Pixel = 194;
			8811: Pixel = 192;
			8812: Pixel = 93;
			8813: Pixel = 29;
			8814: Pixel = 46;
			8815: Pixel = 47;
			8816: Pixel = 51;
			8817: Pixel = 53;
			8818: Pixel = 54;
			8819: Pixel = 54;
			8820: Pixel = 47;
			8821: Pixel = 45;
			8822: Pixel = 51;
			8823: Pixel = 52;
			8824: Pixel = 47;
			8825: Pixel = 83;
			8826: Pixel = 141;
			8827: Pixel = 145;
			8828: Pixel = 142;
			8829: Pixel = 160;
			8830: Pixel = 165;
			8831: Pixel = 165;
			8832: Pixel = 164;
			8833: Pixel = 165;
			8834: Pixel = 164;
			8835: Pixel = 162;
			8836: Pixel = 162;
			8837: Pixel = 161;
			8838: Pixel = 159;
			8839: Pixel = 158;
			8840: Pixel = 158;
			8841: Pixel = 156;
			8842: Pixel = 157;
			8843: Pixel = 157;
			8844: Pixel = 156;
			8845: Pixel = 155;
			8846: Pixel = 154;
			8847: Pixel = 153;
			8848: Pixel = 153;
			8849: Pixel = 152;
			8850: Pixel = 107;
			8851: Pixel = 107;
			8852: Pixel = 106;
			8853: Pixel = 104;
			8854: Pixel = 100;
			8855: Pixel = 99;
			8856: Pixel = 99;
			8857: Pixel = 108;
			8858: Pixel = 128;
			8859: Pixel = 148;
			8860: Pixel = 164;
			8861: Pixel = 171;
			8862: Pixel = 170;
			8863: Pixel = 172;
			8864: Pixel = 172;
			8865: Pixel = 170;
			8866: Pixel = 159;
			8867: Pixel = 142;
			8868: Pixel = 108;
			8869: Pixel = 74;
			8870: Pixel = 73;
			8871: Pixel = 85;
			8872: Pixel = 90;
			8873: Pixel = 93;
			8874: Pixel = 95;
			8875: Pixel = 97;
			8876: Pixel = 97;
			8877: Pixel = 95;
			8878: Pixel = 98;
			8879: Pixel = 97;
			8880: Pixel = 97;
			8881: Pixel = 100;
			8882: Pixel = 104;
			8883: Pixel = 105;
			8884: Pixel = 103;
			8885: Pixel = 90;
			8886: Pixel = 98;
			8887: Pixel = 205;
			8888: Pixel = 213;
			8889: Pixel = 183;
			8890: Pixel = 164;
			8891: Pixel = 185;
			8892: Pixel = 128;
			8893: Pixel = 113;
			8894: Pixel = 136;
			8895: Pixel = 128;
			8896: Pixel = 120;
			8897: Pixel = 110;
			8898: Pixel = 128;
			8899: Pixel = 128;
			8900: Pixel = 122;
			8901: Pixel = 119;
			8902: Pixel = 124;
			8903: Pixel = 135;
			8904: Pixel = 124;
			8905: Pixel = 122;
			8906: Pixel = 101;
			8907: Pixel = 73;
			8908: Pixel = 70;
			8909: Pixel = 69;
			8910: Pixel = 82;
			8911: Pixel = 78;
			8912: Pixel = 59;
			8913: Pixel = 43;
			8914: Pixel = 86;
			8915: Pixel = 78;
			8916: Pixel = 29;
			8917: Pixel = 60;
			8918: Pixel = 90;
			8919: Pixel = 52;
			8920: Pixel = 46;
			8921: Pixel = 64;
			8922: Pixel = 59;
			8923: Pixel = 78;
			8924: Pixel = 61;
			8925: Pixel = 79;
			8926: Pixel = 101;
			8927: Pixel = 66;
			8928: Pixel = 139;
			8929: Pixel = 119;
			8930: Pixel = 167;
			8931: Pixel = 200;
			8932: Pixel = 195;
			8933: Pixel = 189;
			8934: Pixel = 187;
			8935: Pixel = 182;
			8936: Pixel = 180;
			8937: Pixel = 181;
			8938: Pixel = 180;
			8939: Pixel = 170;
			8940: Pixel = 175;
			8941: Pixel = 180;
			8942: Pixel = 180;
			8943: Pixel = 190;
			8944: Pixel = 191;
			8945: Pixel = 187;
			8946: Pixel = 188;
			8947: Pixel = 170;
			8948: Pixel = 89;
			8949: Pixel = 74;
			8950: Pixel = 90;
			8951: Pixel = 95;
			8952: Pixel = 101;
			8953: Pixel = 130;
			8954: Pixel = 113;
			8955: Pixel = 124;
			8956: Pixel = 153;
			8957: Pixel = 164;
			8958: Pixel = 174;
			8959: Pixel = 200;
			8960: Pixel = 167;
			8961: Pixel = 60;
			8962: Pixel = 34;
			8963: Pixel = 42;
			8964: Pixel = 46;
			8965: Pixel = 50;
			8966: Pixel = 52;
			8967: Pixel = 57;
			8968: Pixel = 58;
			8969: Pixel = 50;
			8970: Pixel = 48;
			8971: Pixel = 45;
			8972: Pixel = 52;
			8973: Pixel = 51;
			8974: Pixel = 57;
			8975: Pixel = 107;
			8976: Pixel = 140;
			8977: Pixel = 134;
			8978: Pixel = 146;
			8979: Pixel = 165;
			8980: Pixel = 166;
			8981: Pixel = 165;
			8982: Pixel = 165;
			8983: Pixel = 164;
			8984: Pixel = 161;
			8985: Pixel = 163;
			8986: Pixel = 163;
			8987: Pixel = 162;
			8988: Pixel = 160;
			8989: Pixel = 159;
			8990: Pixel = 158;
			8991: Pixel = 158;
			8992: Pixel = 158;
			8993: Pixel = 157;
			8994: Pixel = 156;
			8995: Pixel = 156;
			8996: Pixel = 155;
			8997: Pixel = 153;
			8998: Pixel = 151;
			8999: Pixel = 151;
			9000: Pixel = 108;
			9001: Pixel = 107;
			9002: Pixel = 106;
			9003: Pixel = 104;
			9004: Pixel = 100;
			9005: Pixel = 99;
			9006: Pixel = 95;
			9007: Pixel = 104;
			9008: Pixel = 127;
			9009: Pixel = 147;
			9010: Pixel = 163;
			9011: Pixel = 170;
			9012: Pixel = 172;
			9013: Pixel = 173;
			9014: Pixel = 173;
			9015: Pixel = 170;
			9016: Pixel = 160;
			9017: Pixel = 141;
			9018: Pixel = 106;
			9019: Pixel = 75;
			9020: Pixel = 75;
			9021: Pixel = 83;
			9022: Pixel = 89;
			9023: Pixel = 93;
			9024: Pixel = 97;
			9025: Pixel = 98;
			9026: Pixel = 97;
			9027: Pixel = 97;
			9028: Pixel = 98;
			9029: Pixel = 97;
			9030: Pixel = 98;
			9031: Pixel = 101;
			9032: Pixel = 105;
			9033: Pixel = 106;
			9034: Pixel = 105;
			9035: Pixel = 103;
			9036: Pixel = 81;
			9037: Pixel = 135;
			9038: Pixel = 219;
			9039: Pixel = 193;
			9040: Pixel = 188;
			9041: Pixel = 175;
			9042: Pixel = 125;
			9043: Pixel = 132;
			9044: Pixel = 124;
			9045: Pixel = 130;
			9046: Pixel = 115;
			9047: Pixel = 123;
			9048: Pixel = 130;
			9049: Pixel = 133;
			9050: Pixel = 127;
			9051: Pixel = 122;
			9052: Pixel = 123;
			9053: Pixel = 126;
			9054: Pixel = 124;
			9055: Pixel = 112;
			9056: Pixel = 96;
			9057: Pixel = 92;
			9058: Pixel = 75;
			9059: Pixel = 80;
			9060: Pixel = 89;
			9061: Pixel = 50;
			9062: Pixel = 37;
			9063: Pixel = 47;
			9064: Pixel = 112;
			9065: Pixel = 58;
			9066: Pixel = 38;
			9067: Pixel = 65;
			9068: Pixel = 76;
			9069: Pixel = 53;
			9070: Pixel = 61;
			9071: Pixel = 60;
			9072: Pixel = 47;
			9073: Pixel = 85;
			9074: Pixel = 61;
			9075: Pixel = 95;
			9076: Pixel = 122;
			9077: Pixel = 124;
			9078: Pixel = 97;
			9079: Pixel = 161;
			9080: Pixel = 200;
			9081: Pixel = 192;
			9082: Pixel = 191;
			9083: Pixel = 186;
			9084: Pixel = 182;
			9085: Pixel = 178;
			9086: Pixel = 179;
			9087: Pixel = 182;
			9088: Pixel = 175;
			9089: Pixel = 169;
			9090: Pixel = 180;
			9091: Pixel = 183;
			9092: Pixel = 183;
			9093: Pixel = 184;
			9094: Pixel = 182;
			9095: Pixel = 184;
			9096: Pixel = 192;
			9097: Pixel = 190;
			9098: Pixel = 138;
			9099: Pixel = 83;
			9100: Pixel = 91;
			9101: Pixel = 108;
			9102: Pixel = 95;
			9103: Pixel = 124;
			9104: Pixel = 127;
			9105: Pixel = 120;
			9106: Pixel = 152;
			9107: Pixel = 182;
			9108: Pixel = 194;
			9109: Pixel = 137;
			9110: Pixel = 48;
			9111: Pixel = 37;
			9112: Pixel = 46;
			9113: Pixel = 46;
			9114: Pixel = 54;
			9115: Pixel = 54;
			9116: Pixel = 50;
			9117: Pixel = 55;
			9118: Pixel = 53;
			9119: Pixel = 46;
			9120: Pixel = 46;
			9121: Pixel = 48;
			9122: Pixel = 55;
			9123: Pixel = 53;
			9124: Pixel = 77;
			9125: Pixel = 126;
			9126: Pixel = 131;
			9127: Pixel = 125;
			9128: Pixel = 156;
			9129: Pixel = 168;
			9130: Pixel = 167;
			9131: Pixel = 164;
			9132: Pixel = 162;
			9133: Pixel = 163;
			9134: Pixel = 161;
			9135: Pixel = 163;
			9136: Pixel = 163;
			9137: Pixel = 162;
			9138: Pixel = 160;
			9139: Pixel = 160;
			9140: Pixel = 159;
			9141: Pixel = 158;
			9142: Pixel = 159;
			9143: Pixel = 159;
			9144: Pixel = 157;
			9145: Pixel = 156;
			9146: Pixel = 155;
			9147: Pixel = 154;
			9148: Pixel = 153;
			9149: Pixel = 152;
			9150: Pixel = 107;
			9151: Pixel = 108;
			9152: Pixel = 104;
			9153: Pixel = 102;
			9154: Pixel = 101;
			9155: Pixel = 99;
			9156: Pixel = 94;
			9157: Pixel = 100;
			9158: Pixel = 125;
			9159: Pixel = 147;
			9160: Pixel = 163;
			9161: Pixel = 171;
			9162: Pixel = 172;
			9163: Pixel = 172;
			9164: Pixel = 175;
			9165: Pixel = 173;
			9166: Pixel = 160;
			9167: Pixel = 142;
			9168: Pixel = 108;
			9169: Pixel = 74;
			9170: Pixel = 71;
			9171: Pixel = 83;
			9172: Pixel = 88;
			9173: Pixel = 93;
			9174: Pixel = 96;
			9175: Pixel = 95;
			9176: Pixel = 96;
			9177: Pixel = 97;
			9178: Pixel = 98;
			9179: Pixel = 99;
			9180: Pixel = 98;
			9181: Pixel = 103;
			9182: Pixel = 106;
			9183: Pixel = 109;
			9184: Pixel = 110;
			9185: Pixel = 106;
			9186: Pixel = 95;
			9187: Pixel = 89;
			9188: Pixel = 194;
			9189: Pixel = 204;
			9190: Pixel = 196;
			9191: Pixel = 171;
			9192: Pixel = 131;
			9193: Pixel = 127;
			9194: Pixel = 116;
			9195: Pixel = 111;
			9196: Pixel = 118;
			9197: Pixel = 132;
			9198: Pixel = 125;
			9199: Pixel = 114;
			9200: Pixel = 117;
			9201: Pixel = 129;
			9202: Pixel = 125;
			9203: Pixel = 121;
			9204: Pixel = 114;
			9205: Pixel = 79;
			9206: Pixel = 68;
			9207: Pixel = 75;
			9208: Pixel = 82;
			9209: Pixel = 98;
			9210: Pixel = 75;
			9211: Pixel = 53;
			9212: Pixel = 45;
			9213: Pixel = 56;
			9214: Pixel = 97;
			9215: Pixel = 51;
			9216: Pixel = 64;
			9217: Pixel = 61;
			9218: Pixel = 46;
			9219: Pixel = 54;
			9220: Pixel = 67;
			9221: Pixel = 76;
			9222: Pixel = 67;
			9223: Pixel = 83;
			9224: Pixel = 72;
			9225: Pixel = 94;
			9226: Pixel = 116;
			9227: Pixel = 124;
			9228: Pixel = 149;
			9229: Pixel = 182;
			9230: Pixel = 184;
			9231: Pixel = 183;
			9232: Pixel = 187;
			9233: Pixel = 180;
			9234: Pixel = 174;
			9235: Pixel = 176;
			9236: Pixel = 175;
			9237: Pixel = 174;
			9238: Pixel = 174;
			9239: Pixel = 175;
			9240: Pixel = 179;
			9241: Pixel = 180;
			9242: Pixel = 184;
			9243: Pixel = 188;
			9244: Pixel = 190;
			9245: Pixel = 194;
			9246: Pixel = 199;
			9247: Pixel = 196;
			9248: Pixel = 168;
			9249: Pixel = 109;
			9250: Pixel = 78;
			9251: Pixel = 97;
			9252: Pixel = 101;
			9253: Pixel = 84;
			9254: Pixel = 133;
			9255: Pixel = 132;
			9256: Pixel = 151;
			9257: Pixel = 168;
			9258: Pixel = 105;
			9259: Pixel = 34;
			9260: Pixel = 42;
			9261: Pixel = 48;
			9262: Pixel = 45;
			9263: Pixel = 49;
			9264: Pixel = 57;
			9265: Pixel = 55;
			9266: Pixel = 55;
			9267: Pixel = 56;
			9268: Pixel = 51;
			9269: Pixel = 43;
			9270: Pixel = 48;
			9271: Pixel = 52;
			9272: Pixel = 50;
			9273: Pixel = 57;
			9274: Pixel = 97;
			9275: Pixel = 134;
			9276: Pixel = 124;
			9277: Pixel = 133;
			9278: Pixel = 164;
			9279: Pixel = 168;
			9280: Pixel = 166;
			9281: Pixel = 163;
			9282: Pixel = 163;
			9283: Pixel = 163;
			9284: Pixel = 163;
			9285: Pixel = 163;
			9286: Pixel = 160;
			9287: Pixel = 161;
			9288: Pixel = 162;
			9289: Pixel = 160;
			9290: Pixel = 159;
			9291: Pixel = 159;
			9292: Pixel = 159;
			9293: Pixel = 157;
			9294: Pixel = 157;
			9295: Pixel = 156;
			9296: Pixel = 155;
			9297: Pixel = 154;
			9298: Pixel = 153;
			9299: Pixel = 151;
			9300: Pixel = 107;
			9301: Pixel = 107;
			9302: Pixel = 104;
			9303: Pixel = 103;
			9304: Pixel = 101;
			9305: Pixel = 99;
			9306: Pixel = 92;
			9307: Pixel = 97;
			9308: Pixel = 124;
			9309: Pixel = 147;
			9310: Pixel = 160;
			9311: Pixel = 170;
			9312: Pixel = 172;
			9313: Pixel = 172;
			9314: Pixel = 174;
			9315: Pixel = 172;
			9316: Pixel = 162;
			9317: Pixel = 142;
			9318: Pixel = 110;
			9319: Pixel = 73;
			9320: Pixel = 72;
			9321: Pixel = 81;
			9322: Pixel = 88;
			9323: Pixel = 92;
			9324: Pixel = 97;
			9325: Pixel = 97;
			9326: Pixel = 97;
			9327: Pixel = 95;
			9328: Pixel = 96;
			9329: Pixel = 97;
			9330: Pixel = 99;
			9331: Pixel = 102;
			9332: Pixel = 105;
			9333: Pixel = 110;
			9334: Pixel = 112;
			9335: Pixel = 108;
			9336: Pixel = 103;
			9337: Pixel = 83;
			9338: Pixel = 176;
			9339: Pixel = 221;
			9340: Pixel = 199;
			9341: Pixel = 188;
			9342: Pixel = 136;
			9343: Pixel = 122;
			9344: Pixel = 118;
			9345: Pixel = 105;
			9346: Pixel = 124;
			9347: Pixel = 124;
			9348: Pixel = 115;
			9349: Pixel = 120;
			9350: Pixel = 133;
			9351: Pixel = 131;
			9352: Pixel = 109;
			9353: Pixel = 128;
			9354: Pixel = 106;
			9355: Pixel = 68;
			9356: Pixel = 66;
			9357: Pixel = 56;
			9358: Pixel = 66;
			9359: Pixel = 86;
			9360: Pixel = 70;
			9361: Pixel = 60;
			9362: Pixel = 51;
			9363: Pixel = 64;
			9364: Pixel = 72;
			9365: Pixel = 95;
			9366: Pixel = 61;
			9367: Pixel = 44;
			9368: Pixel = 48;
			9369: Pixel = 47;
			9370: Pixel = 49;
			9371: Pixel = 47;
			9372: Pixel = 38;
			9373: Pixel = 61;
			9374: Pixel = 94;
			9375: Pixel = 77;
			9376: Pixel = 97;
			9377: Pixel = 136;
			9378: Pixel = 157;
			9379: Pixel = 175;
			9380: Pixel = 176;
			9381: Pixel = 181;
			9382: Pixel = 179;
			9383: Pixel = 170;
			9384: Pixel = 168;
			9385: Pixel = 175;
			9386: Pixel = 173;
			9387: Pixel = 176;
			9388: Pixel = 175;
			9389: Pixel = 172;
			9390: Pixel = 170;
			9391: Pixel = 185;
			9392: Pixel = 197;
			9393: Pixel = 195;
			9394: Pixel = 195;
			9395: Pixel = 197;
			9396: Pixel = 196;
			9397: Pixel = 199;
			9398: Pixel = 186;
			9399: Pixel = 132;
			9400: Pixel = 88;
			9401: Pixel = 58;
			9402: Pixel = 81;
			9403: Pixel = 83;
			9404: Pixel = 100;
			9405: Pixel = 138;
			9406: Pixel = 149;
			9407: Pixel = 135;
			9408: Pixel = 78;
			9409: Pixel = 39;
			9410: Pixel = 43;
			9411: Pixel = 42;
			9412: Pixel = 50;
			9413: Pixel = 55;
			9414: Pixel = 54;
			9415: Pixel = 58;
			9416: Pixel = 58;
			9417: Pixel = 55;
			9418: Pixel = 48;
			9419: Pixel = 41;
			9420: Pixel = 49;
			9421: Pixel = 52;
			9422: Pixel = 50;
			9423: Pixel = 70;
			9424: Pixel = 121;
			9425: Pixel = 133;
			9426: Pixel = 121;
			9427: Pixel = 142;
			9428: Pixel = 165;
			9429: Pixel = 166;
			9430: Pixel = 166;
			9431: Pixel = 165;
			9432: Pixel = 165;
			9433: Pixel = 162;
			9434: Pixel = 163;
			9435: Pixel = 164;
			9436: Pixel = 162;
			9437: Pixel = 162;
			9438: Pixel = 162;
			9439: Pixel = 160;
			9440: Pixel = 161;
			9441: Pixel = 162;
			9442: Pixel = 159;
			9443: Pixel = 157;
			9444: Pixel = 157;
			9445: Pixel = 157;
			9446: Pixel = 156;
			9447: Pixel = 154;
			9448: Pixel = 153;
			9449: Pixel = 152;
			9450: Pixel = 106;
			9451: Pixel = 104;
			9452: Pixel = 105;
			9453: Pixel = 104;
			9454: Pixel = 99;
			9455: Pixel = 98;
			9456: Pixel = 90;
			9457: Pixel = 96;
			9458: Pixel = 123;
			9459: Pixel = 145;
			9460: Pixel = 160;
			9461: Pixel = 170;
			9462: Pixel = 171;
			9463: Pixel = 173;
			9464: Pixel = 174;
			9465: Pixel = 173;
			9466: Pixel = 161;
			9467: Pixel = 143;
			9468: Pixel = 109;
			9469: Pixel = 74;
			9470: Pixel = 73;
			9471: Pixel = 84;
			9472: Pixel = 91;
			9473: Pixel = 94;
			9474: Pixel = 98;
			9475: Pixel = 99;
			9476: Pixel = 100;
			9477: Pixel = 98;
			9478: Pixel = 99;
			9479: Pixel = 97;
			9480: Pixel = 98;
			9481: Pixel = 103;
			9482: Pixel = 106;
			9483: Pixel = 113;
			9484: Pixel = 113;
			9485: Pixel = 110;
			9486: Pixel = 104;
			9487: Pixel = 85;
			9488: Pixel = 175;
			9489: Pixel = 221;
			9490: Pixel = 212;
			9491: Pixel = 162;
			9492: Pixel = 108;
			9493: Pixel = 124;
			9494: Pixel = 118;
			9495: Pixel = 124;
			9496: Pixel = 117;
			9497: Pixel = 107;
			9498: Pixel = 130;
			9499: Pixel = 138;
			9500: Pixel = 131;
			9501: Pixel = 123;
			9502: Pixel = 91;
			9503: Pixel = 83;
			9504: Pixel = 68;
			9505: Pixel = 81;
			9506: Pixel = 55;
			9507: Pixel = 45;
			9508: Pixel = 49;
			9509: Pixel = 77;
			9510: Pixel = 71;
			9511: Pixel = 84;
			9512: Pixel = 56;
			9513: Pixel = 63;
			9514: Pixel = 54;
			9515: Pixel = 118;
			9516: Pixel = 82;
			9517: Pixel = 37;
			9518: Pixel = 47;
			9519: Pixel = 47;
			9520: Pixel = 47;
			9521: Pixel = 39;
			9522: Pixel = 40;
			9523: Pixel = 101;
			9524: Pixel = 99;
			9525: Pixel = 99;
			9526: Pixel = 141;
			9527: Pixel = 166;
			9528: Pixel = 179;
			9529: Pixel = 179;
			9530: Pixel = 185;
			9531: Pixel = 186;
			9532: Pixel = 172;
			9533: Pixel = 163;
			9534: Pixel = 168;
			9535: Pixel = 175;
			9536: Pixel = 180;
			9537: Pixel = 164;
			9538: Pixel = 166;
			9539: Pixel = 173;
			9540: Pixel = 186;
			9541: Pixel = 196;
			9542: Pixel = 199;
			9543: Pixel = 197;
			9544: Pixel = 195;
			9545: Pixel = 197;
			9546: Pixel = 198;
			9547: Pixel = 198;
			9548: Pixel = 187;
			9549: Pixel = 146;
			9550: Pixel = 96;
			9551: Pixel = 64;
			9552: Pixel = 45;
			9553: Pixel = 83;
			9554: Pixel = 85;
			9555: Pixel = 130;
			9556: Pixel = 147;
			9557: Pixel = 143;
			9558: Pixel = 69;
			9559: Pixel = 43;
			9560: Pixel = 44;
			9561: Pixel = 46;
			9562: Pixel = 49;
			9563: Pixel = 57;
			9564: Pixel = 56;
			9565: Pixel = 58;
			9566: Pixel = 61;
			9567: Pixel = 53;
			9568: Pixel = 48;
			9569: Pixel = 43;
			9570: Pixel = 48;
			9571: Pixel = 49;
			9572: Pixel = 47;
			9573: Pixel = 91;
			9574: Pixel = 136;
			9575: Pixel = 129;
			9576: Pixel = 127;
			9577: Pixel = 153;
			9578: Pixel = 161;
			9579: Pixel = 165;
			9580: Pixel = 165;
			9581: Pixel = 164;
			9582: Pixel = 164;
			9583: Pixel = 162;
			9584: Pixel = 160;
			9585: Pixel = 162;
			9586: Pixel = 162;
			9587: Pixel = 163;
			9588: Pixel = 162;
			9589: Pixel = 161;
			9590: Pixel = 160;
			9591: Pixel = 159;
			9592: Pixel = 159;
			9593: Pixel = 158;
			9594: Pixel = 159;
			9595: Pixel = 158;
			9596: Pixel = 157;
			9597: Pixel = 155;
			9598: Pixel = 152;
			9599: Pixel = 151;
			9600: Pixel = 105;
			9601: Pixel = 105;
			9602: Pixel = 105;
			9603: Pixel = 104;
			9604: Pixel = 100;
			9605: Pixel = 98;
			9606: Pixel = 91;
			9607: Pixel = 95;
			9608: Pixel = 123;
			9609: Pixel = 145;
			9610: Pixel = 161;
			9611: Pixel = 169;
			9612: Pixel = 172;
			9613: Pixel = 174;
			9614: Pixel = 173;
			9615: Pixel = 171;
			9616: Pixel = 160;
			9617: Pixel = 143;
			9618: Pixel = 109;
			9619: Pixel = 77;
			9620: Pixel = 73;
			9621: Pixel = 83;
			9622: Pixel = 93;
			9623: Pixel = 96;
			9624: Pixel = 98;
			9625: Pixel = 99;
			9626: Pixel = 100;
			9627: Pixel = 100;
			9628: Pixel = 98;
			9629: Pixel = 99;
			9630: Pixel = 100;
			9631: Pixel = 105;
			9632: Pixel = 107;
			9633: Pixel = 111;
			9634: Pixel = 114;
			9635: Pixel = 112;
			9636: Pixel = 108;
			9637: Pixel = 88;
			9638: Pixel = 167;
			9639: Pixel = 224;
			9640: Pixel = 206;
			9641: Pixel = 121;
			9642: Pixel = 100;
			9643: Pixel = 115;
			9644: Pixel = 117;
			9645: Pixel = 119;
			9646: Pixel = 110;
			9647: Pixel = 125;
			9648: Pixel = 129;
			9649: Pixel = 130;
			9650: Pixel = 122;
			9651: Pixel = 128;
			9652: Pixel = 74;
			9653: Pixel = 37;
			9654: Pixel = 66;
			9655: Pixel = 66;
			9656: Pixel = 42;
			9657: Pixel = 46;
			9658: Pixel = 45;
			9659: Pixel = 70;
			9660: Pixel = 75;
			9661: Pixel = 78;
			9662: Pixel = 61;
			9663: Pixel = 66;
			9664: Pixel = 47;
			9665: Pixel = 74;
			9666: Pixel = 123;
			9667: Pixel = 77;
			9668: Pixel = 63;
			9669: Pixel = 40;
			9670: Pixel = 36;
			9671: Pixel = 32;
			9672: Pixel = 114;
			9673: Pixel = 114;
			9674: Pixel = 113;
			9675: Pixel = 163;
			9676: Pixel = 140;
			9677: Pixel = 179;
			9678: Pixel = 181;
			9679: Pixel = 187;
			9680: Pixel = 192;
			9681: Pixel = 178;
			9682: Pixel = 164;
			9683: Pixel = 159;
			9684: Pixel = 167;
			9685: Pixel = 182;
			9686: Pixel = 172;
			9687: Pixel = 159;
			9688: Pixel = 171;
			9689: Pixel = 184;
			9690: Pixel = 192;
			9691: Pixel = 195;
			9692: Pixel = 199;
			9693: Pixel = 201;
			9694: Pixel = 199;
			9695: Pixel = 200;
			9696: Pixel = 203;
			9697: Pixel = 203;
			9698: Pixel = 196;
			9699: Pixel = 157;
			9700: Pixel = 102;
			9701: Pixel = 67;
			9702: Pixel = 39;
			9703: Pixel = 62;
			9704: Pixel = 76;
			9705: Pixel = 125;
			9706: Pixel = 159;
			9707: Pixel = 136;
			9708: Pixel = 51;
			9709: Pixel = 46;
			9710: Pixel = 46;
			9711: Pixel = 47;
			9712: Pixel = 50;
			9713: Pixel = 55;
			9714: Pixel = 58;
			9715: Pixel = 62;
			9716: Pixel = 61;
			9717: Pixel = 51;
			9718: Pixel = 44;
			9719: Pixel = 45;
			9720: Pixel = 51;
			9721: Pixel = 46;
			9722: Pixel = 58;
			9723: Pixel = 116;
			9724: Pixel = 141;
			9725: Pixel = 128;
			9726: Pixel = 141;
			9727: Pixel = 153;
			9728: Pixel = 151;
			9729: Pixel = 159;
			9730: Pixel = 164;
			9731: Pixel = 164;
			9732: Pixel = 166;
			9733: Pixel = 164;
			9734: Pixel = 161;
			9735: Pixel = 161;
			9736: Pixel = 161;
			9737: Pixel = 162;
			9738: Pixel = 163;
			9739: Pixel = 162;
			9740: Pixel = 160;
			9741: Pixel = 159;
			9742: Pixel = 158;
			9743: Pixel = 157;
			9744: Pixel = 158;
			9745: Pixel = 157;
			9746: Pixel = 157;
			9747: Pixel = 155;
			9748: Pixel = 154;
			9749: Pixel = 150;
			9750: Pixel = 102;
			9751: Pixel = 104;
			9752: Pixel = 103;
			9753: Pixel = 101;
			9754: Pixel = 100;
			9755: Pixel = 100;
			9756: Pixel = 93;
			9757: Pixel = 97;
			9758: Pixel = 124;
			9759: Pixel = 145;
			9760: Pixel = 160;
			9761: Pixel = 170;
			9762: Pixel = 172;
			9763: Pixel = 172;
			9764: Pixel = 174;
			9765: Pixel = 172;
			9766: Pixel = 162;
			9767: Pixel = 145;
			9768: Pixel = 113;
			9769: Pixel = 77;
			9770: Pixel = 74;
			9771: Pixel = 82;
			9772: Pixel = 91;
			9773: Pixel = 94;
			9774: Pixel = 99;
			9775: Pixel = 99;
			9776: Pixel = 101;
			9777: Pixel = 101;
			9778: Pixel = 99;
			9779: Pixel = 100;
			9780: Pixel = 103;
			9781: Pixel = 102;
			9782: Pixel = 106;
			9783: Pixel = 116;
			9784: Pixel = 115;
			9785: Pixel = 114;
			9786: Pixel = 112;
			9787: Pixel = 94;
			9788: Pixel = 135;
			9789: Pixel = 229;
			9790: Pixel = 185;
			9791: Pixel = 105;
			9792: Pixel = 110;
			9793: Pixel = 110;
			9794: Pixel = 111;
			9795: Pixel = 113;
			9796: Pixel = 128;
			9797: Pixel = 127;
			9798: Pixel = 111;
			9799: Pixel = 95;
			9800: Pixel = 102;
			9801: Pixel = 94;
			9802: Pixel = 75;
			9803: Pixel = 48;
			9804: Pixel = 87;
			9805: Pixel = 46;
			9806: Pixel = 42;
			9807: Pixel = 51;
			9808: Pixel = 50;
			9809: Pixel = 47;
			9810: Pixel = 70;
			9811: Pixel = 70;
			9812: Pixel = 64;
			9813: Pixel = 76;
			9814: Pixel = 55;
			9815: Pixel = 54;
			9816: Pixel = 115;
			9817: Pixel = 60;
			9818: Pixel = 52;
			9819: Pixel = 36;
			9820: Pixel = 25;
			9821: Pixel = 108;
			9822: Pixel = 138;
			9823: Pixel = 125;
			9824: Pixel = 176;
			9825: Pixel = 165;
			9826: Pixel = 134;
			9827: Pixel = 165;
			9828: Pixel = 174;
			9829: Pixel = 187;
			9830: Pixel = 182;
			9831: Pixel = 170;
			9832: Pixel = 164;
			9833: Pixel = 162;
			9834: Pixel = 177;
			9835: Pixel = 170;
			9836: Pixel = 157;
			9837: Pixel = 169;
			9838: Pixel = 179;
			9839: Pixel = 187;
			9840: Pixel = 195;
			9841: Pixel = 196;
			9842: Pixel = 200;
			9843: Pixel = 201;
			9844: Pixel = 201;
			9845: Pixel = 205;
			9846: Pixel = 209;
			9847: Pixel = 209;
			9848: Pixel = 205;
			9849: Pixel = 175;
			9850: Pixel = 117;
			9851: Pixel = 76;
			9852: Pixel = 40;
			9853: Pixel = 49;
			9854: Pixel = 67;
			9855: Pixel = 108;
			9856: Pixel = 171;
			9857: Pixel = 132;
			9858: Pixel = 47;
			9859: Pixel = 47;
			9860: Pixel = 50;
			9861: Pixel = 52;
			9862: Pixel = 53;
			9863: Pixel = 54;
			9864: Pixel = 57;
			9865: Pixel = 62;
			9866: Pixel = 57;
			9867: Pixel = 45;
			9868: Pixel = 45;
			9869: Pixel = 50;
			9870: Pixel = 50;
			9871: Pixel = 45;
			9872: Pixel = 81;
			9873: Pixel = 138;
			9874: Pixel = 135;
			9875: Pixel = 132;
			9876: Pixel = 155;
			9877: Pixel = 153;
			9878: Pixel = 150;
			9879: Pixel = 150;
			9880: Pixel = 153;
			9881: Pixel = 157;
			9882: Pixel = 160;
			9883: Pixel = 160;
			9884: Pixel = 161;
			9885: Pixel = 162;
			9886: Pixel = 160;
			9887: Pixel = 160;
			9888: Pixel = 162;
			9889: Pixel = 163;
			9890: Pixel = 159;
			9891: Pixel = 159;
			9892: Pixel = 159;
			9893: Pixel = 157;
			9894: Pixel = 157;
			9895: Pixel = 157;
			9896: Pixel = 156;
			9897: Pixel = 155;
			9898: Pixel = 153;
			9899: Pixel = 150;
			9900: Pixel = 103;
			9901: Pixel = 104;
			9902: Pixel = 103;
			9903: Pixel = 103;
			9904: Pixel = 100;
			9905: Pixel = 98;
			9906: Pixel = 93;
			9907: Pixel = 95;
			9908: Pixel = 123;
			9909: Pixel = 146;
			9910: Pixel = 161;
			9911: Pixel = 169;
			9912: Pixel = 172;
			9913: Pixel = 173;
			9914: Pixel = 174;
			9915: Pixel = 173;
			9916: Pixel = 163;
			9917: Pixel = 142;
			9918: Pixel = 113;
			9919: Pixel = 80;
			9920: Pixel = 74;
			9921: Pixel = 82;
			9922: Pixel = 90;
			9923: Pixel = 95;
			9924: Pixel = 101;
			9925: Pixel = 102;
			9926: Pixel = 104;
			9927: Pixel = 103;
			9928: Pixel = 101;
			9929: Pixel = 100;
			9930: Pixel = 99;
			9931: Pixel = 99;
			9932: Pixel = 136;
			9933: Pixel = 127;
			9934: Pixel = 111;
			9935: Pixel = 115;
			9936: Pixel = 114;
			9937: Pixel = 106;
			9938: Pixel = 107;
			9939: Pixel = 214;
			9940: Pixel = 176;
			9941: Pixel = 105;
			9942: Pixel = 121;
			9943: Pixel = 115;
			9944: Pixel = 104;
			9945: Pixel = 125;
			9946: Pixel = 131;
			9947: Pixel = 125;
			9948: Pixel = 102;
			9949: Pixel = 83;
			9950: Pixel = 73;
			9951: Pixel = 55;
			9952: Pixel = 58;
			9953: Pixel = 60;
			9954: Pixel = 84;
			9955: Pixel = 37;
			9956: Pixel = 56;
			9957: Pixel = 61;
			9958: Pixel = 50;
			9959: Pixel = 49;
			9960: Pixel = 51;
			9961: Pixel = 60;
			9962: Pixel = 55;
			9963: Pixel = 79;
			9964: Pixel = 97;
			9965: Pixel = 54;
			9966: Pixel = 93;
			9967: Pixel = 59;
			9968: Pixel = 30;
			9969: Pixel = 27;
			9970: Pixel = 92;
			9971: Pixel = 145;
			9972: Pixel = 122;
			9973: Pixel = 177;
			9974: Pixel = 171;
			9975: Pixel = 164;
			9976: Pixel = 147;
			9977: Pixel = 164;
			9978: Pixel = 172;
			9979: Pixel = 189;
			9980: Pixel = 178;
			9981: Pixel = 169;
			9982: Pixel = 171;
			9983: Pixel = 171;
			9984: Pixel = 159;
			9985: Pixel = 152;
			9986: Pixel = 166;
			9987: Pixel = 173;
			9988: Pixel = 184;
			9989: Pixel = 189;
			9990: Pixel = 195;
			9991: Pixel = 198;
			9992: Pixel = 200;
			9993: Pixel = 201;
			9994: Pixel = 202;
			9995: Pixel = 207;
			9996: Pixel = 208;
			9997: Pixel = 211;
			9998: Pixel = 208;
			9999: Pixel = 188;
			10000: Pixel = 134;
			10001: Pixel = 84;
			10002: Pixel = 49;
			10003: Pixel = 38;
			10004: Pixel = 54;
			10005: Pixel = 81;
			10006: Pixel = 161;
			10007: Pixel = 146;
			10008: Pixel = 58;
			10009: Pixel = 52;
			10010: Pixel = 50;
			10011: Pixel = 53;
			10012: Pixel = 56;
			10013: Pixel = 57;
			10014: Pixel = 61;
			10015: Pixel = 64;
			10016: Pixel = 54;
			10017: Pixel = 45;
			10018: Pixel = 47;
			10019: Pixel = 55;
			10020: Pixel = 49;
			10021: Pixel = 42;
			10022: Pixel = 101;
			10023: Pixel = 144;
			10024: Pixel = 131;
			10025: Pixel = 144;
			10026: Pixel = 162;
			10027: Pixel = 155;
			10028: Pixel = 152;
			10029: Pixel = 151;
			10030: Pixel = 149;
			10031: Pixel = 150;
			10032: Pixel = 149;
			10033: Pixel = 152;
			10034: Pixel = 154;
			10035: Pixel = 158;
			10036: Pixel = 158;
			10037: Pixel = 160;
			10038: Pixel = 160;
			10039: Pixel = 161;
			10040: Pixel = 161;
			10041: Pixel = 160;
			10042: Pixel = 159;
			10043: Pixel = 158;
			10044: Pixel = 156;
			10045: Pixel = 156;
			10046: Pixel = 155;
			10047: Pixel = 155;
			10048: Pixel = 154;
			10049: Pixel = 150;
			10050: Pixel = 106;
			10051: Pixel = 106;
			10052: Pixel = 102;
			10053: Pixel = 99;
			10054: Pixel = 100;
			10055: Pixel = 98;
			10056: Pixel = 92;
			10057: Pixel = 98;
			10058: Pixel = 121;
			10059: Pixel = 144;
			10060: Pixel = 160;
			10061: Pixel = 170;
			10062: Pixel = 173;
			10063: Pixel = 174;
			10064: Pixel = 174;
			10065: Pixel = 174;
			10066: Pixel = 162;
			10067: Pixel = 143;
			10068: Pixel = 113;
			10069: Pixel = 81;
			10070: Pixel = 78;
			10071: Pixel = 86;
			10072: Pixel = 93;
			10073: Pixel = 100;
			10074: Pixel = 101;
			10075: Pixel = 102;
			10076: Pixel = 103;
			10077: Pixel = 102;
			10078: Pixel = 100;
			10079: Pixel = 99;
			10080: Pixel = 100;
			10081: Pixel = 109;
			10082: Pixel = 123;
			10083: Pixel = 111;
			10084: Pixel = 116;
			10085: Pixel = 116;
			10086: Pixel = 116;
			10087: Pixel = 117;
			10088: Pixel = 100;
			10089: Pixel = 164;
			10090: Pixel = 197;
			10091: Pixel = 112;
			10092: Pixel = 112;
			10093: Pixel = 114;
			10094: Pixel = 125;
			10095: Pixel = 123;
			10096: Pixel = 129;
			10097: Pixel = 128;
			10098: Pixel = 111;
			10099: Pixel = 84;
			10100: Pixel = 55;
			10101: Pixel = 56;
			10102: Pixel = 37;
			10103: Pixel = 55;
			10104: Pixel = 77;
			10105: Pixel = 45;
			10106: Pixel = 59;
			10107: Pixel = 56;
			10108: Pixel = 49;
			10109: Pixel = 55;
			10110: Pixel = 50;
			10111: Pixel = 57;
			10112: Pixel = 48;
			10113: Pixel = 80;
			10114: Pixel = 101;
			10115: Pixel = 77;
			10116: Pixel = 100;
			10117: Pixel = 94;
			10118: Pixel = 15;
			10119: Pixel = 79;
			10120: Pixel = 145;
			10121: Pixel = 124;
			10122: Pixel = 173;
			10123: Pixel = 178;
			10124: Pixel = 179;
			10125: Pixel = 175;
			10126: Pixel = 153;
			10127: Pixel = 161;
			10128: Pixel = 179;
			10129: Pixel = 198;
			10130: Pixel = 176;
			10131: Pixel = 167;
			10132: Pixel = 166;
			10133: Pixel = 154;
			10134: Pixel = 152;
			10135: Pixel = 164;
			10136: Pixel = 169;
			10137: Pixel = 175;
			10138: Pixel = 188;
			10139: Pixel = 192;
			10140: Pixel = 195;
			10141: Pixel = 198;
			10142: Pixel = 201;
			10143: Pixel = 203;
			10144: Pixel = 203;
			10145: Pixel = 208;
			10146: Pixel = 209;
			10147: Pixel = 211;
			10148: Pixel = 209;
			10149: Pixel = 197;
			10150: Pixel = 146;
			10151: Pixel = 91;
			10152: Pixel = 54;
			10153: Pixel = 33;
			10154: Pixel = 47;
			10155: Pixel = 73;
			10156: Pixel = 154;
			10157: Pixel = 149;
			10158: Pixel = 66;
			10159: Pixel = 51;
			10160: Pixel = 54;
			10161: Pixel = 54;
			10162: Pixel = 56;
			10163: Pixel = 60;
			10164: Pixel = 62;
			10165: Pixel = 64;
			10166: Pixel = 50;
			10167: Pixel = 45;
			10168: Pixel = 48;
			10169: Pixel = 54;
			10170: Pixel = 43;
			10171: Pixel = 61;
			10172: Pixel = 127;
			10173: Pixel = 142;
			10174: Pixel = 132;
			10175: Pixel = 156;
			10176: Pixel = 165;
			10177: Pixel = 160;
			10178: Pixel = 156;
			10179: Pixel = 154;
			10180: Pixel = 151;
			10181: Pixel = 150;
			10182: Pixel = 148;
			10183: Pixel = 148;
			10184: Pixel = 150;
			10185: Pixel = 149;
			10186: Pixel = 147;
			10187: Pixel = 151;
			10188: Pixel = 154;
			10189: Pixel = 159;
			10190: Pixel = 160;
			10191: Pixel = 159;
			10192: Pixel = 157;
			10193: Pixel = 156;
			10194: Pixel = 155;
			10195: Pixel = 154;
			10196: Pixel = 154;
			10197: Pixel = 153;
			10198: Pixel = 151;
			10199: Pixel = 149;
			10200: Pixel = 104;
			10201: Pixel = 104;
			10202: Pixel = 101;
			10203: Pixel = 99;
			10204: Pixel = 98;
			10205: Pixel = 94;
			10206: Pixel = 90;
			10207: Pixel = 94;
			10208: Pixel = 120;
			10209: Pixel = 143;
			10210: Pixel = 160;
			10211: Pixel = 170;
			10212: Pixel = 173;
			10213: Pixel = 175;
			10214: Pixel = 174;
			10215: Pixel = 172;
			10216: Pixel = 161;
			10217: Pixel = 143;
			10218: Pixel = 112;
			10219: Pixel = 80;
			10220: Pixel = 79;
			10221: Pixel = 90;
			10222: Pixel = 95;
			10223: Pixel = 96;
			10224: Pixel = 100;
			10225: Pixel = 101;
			10226: Pixel = 101;
			10227: Pixel = 103;
			10228: Pixel = 102;
			10229: Pixel = 102;
			10230: Pixel = 103;
			10231: Pixel = 106;
			10232: Pixel = 119;
			10233: Pixel = 113;
			10234: Pixel = 118;
			10235: Pixel = 121;
			10236: Pixel = 120;
			10237: Pixel = 121;
			10238: Pixel = 112;
			10239: Pixel = 125;
			10240: Pixel = 189;
			10241: Pixel = 126;
			10242: Pixel = 109;
			10243: Pixel = 127;
			10244: Pixel = 130;
			10245: Pixel = 131;
			10246: Pixel = 131;
			10247: Pixel = 104;
			10248: Pixel = 69;
			10249: Pixel = 48;
			10250: Pixel = 76;
			10251: Pixel = 66;
			10252: Pixel = 37;
			10253: Pixel = 43;
			10254: Pixel = 82;
			10255: Pixel = 62;
			10256: Pixel = 50;
			10257: Pixel = 65;
			10258: Pixel = 49;
			10259: Pixel = 51;
			10260: Pixel = 56;
			10261: Pixel = 65;
			10262: Pixel = 44;
			10263: Pixel = 72;
			10264: Pixel = 69;
			10265: Pixel = 51;
			10266: Pixel = 66;
			10267: Pixel = 99;
			10268: Pixel = 56;
			10269: Pixel = 143;
			10270: Pixel = 121;
			10271: Pixel = 159;
			10272: Pixel = 172;
			10273: Pixel = 178;
			10274: Pixel = 188;
			10275: Pixel = 183;
			10276: Pixel = 146;
			10277: Pixel = 153;
			10278: Pixel = 188;
			10279: Pixel = 189;
			10280: Pixel = 163;
			10281: Pixel = 160;
			10282: Pixel = 156;
			10283: Pixel = 156;
			10284: Pixel = 164;
			10285: Pixel = 171;
			10286: Pixel = 172;
			10287: Pixel = 177;
			10288: Pixel = 185;
			10289: Pixel = 193;
			10290: Pixel = 195;
			10291: Pixel = 198;
			10292: Pixel = 201;
			10293: Pixel = 203;
			10294: Pixel = 204;
			10295: Pixel = 207;
			10296: Pixel = 209;
			10297: Pixel = 212;
			10298: Pixel = 213;
			10299: Pixel = 204;
			10300: Pixel = 160;
			10301: Pixel = 105;
			10302: Pixel = 66;
			10303: Pixel = 42;
			10304: Pixel = 42;
			10305: Pixel = 60;
			10306: Pixel = 137;
			10307: Pixel = 158;
			10308: Pixel = 72;
			10309: Pixel = 44;
			10310: Pixel = 54;
			10311: Pixel = 57;
			10312: Pixel = 58;
			10313: Pixel = 57;
			10314: Pixel = 60;
			10315: Pixel = 60;
			10316: Pixel = 51;
			10317: Pixel = 46;
			10318: Pixel = 53;
			10319: Pixel = 53;
			10320: Pixel = 41;
			10321: Pixel = 87;
			10322: Pixel = 147;
			10323: Pixel = 136;
			10324: Pixel = 139;
			10325: Pixel = 162;
			10326: Pixel = 165;
			10327: Pixel = 163;
			10328: Pixel = 162;
			10329: Pixel = 158;
			10330: Pixel = 156;
			10331: Pixel = 155;
			10332: Pixel = 153;
			10333: Pixel = 152;
			10334: Pixel = 152;
			10335: Pixel = 148;
			10336: Pixel = 145;
			10337: Pixel = 145;
			10338: Pixel = 144;
			10339: Pixel = 148;
			10340: Pixel = 149;
			10341: Pixel = 152;
			10342: Pixel = 153;
			10343: Pixel = 153;
			10344: Pixel = 153;
			10345: Pixel = 152;
			10346: Pixel = 153;
			10347: Pixel = 154;
			10348: Pixel = 152;
			10349: Pixel = 150;
			10350: Pixel = 102;
			10351: Pixel = 102;
			10352: Pixel = 101;
			10353: Pixel = 100;
			10354: Pixel = 97;
			10355: Pixel = 97;
			10356: Pixel = 90;
			10357: Pixel = 93;
			10358: Pixel = 122;
			10359: Pixel = 144;
			10360: Pixel = 160;
			10361: Pixel = 171;
			10362: Pixel = 173;
			10363: Pixel = 174;
			10364: Pixel = 175;
			10365: Pixel = 172;
			10366: Pixel = 162;
			10367: Pixel = 145;
			10368: Pixel = 110;
			10369: Pixel = 79;
			10370: Pixel = 78;
			10371: Pixel = 88;
			10372: Pixel = 94;
			10373: Pixel = 97;
			10374: Pixel = 101;
			10375: Pixel = 102;
			10376: Pixel = 103;
			10377: Pixel = 105;
			10378: Pixel = 103;
			10379: Pixel = 101;
			10380: Pixel = 104;
			10381: Pixel = 107;
			10382: Pixel = 114;
			10383: Pixel = 116;
			10384: Pixel = 115;
			10385: Pixel = 115;
			10386: Pixel = 114;
			10387: Pixel = 112;
			10388: Pixel = 118;
			10389: Pixel = 122;
			10390: Pixel = 118;
			10391: Pixel = 112;
			10392: Pixel = 122;
			10393: Pixel = 137;
			10394: Pixel = 133;
			10395: Pixel = 127;
			10396: Pixel = 115;
			10397: Pixel = 67;
			10398: Pixel = 58;
			10399: Pixel = 43;
			10400: Pixel = 72;
			10401: Pixel = 61;
			10402: Pixel = 55;
			10403: Pixel = 44;
			10404: Pixel = 47;
			10405: Pixel = 63;
			10406: Pixel = 79;
			10407: Pixel = 58;
			10408: Pixel = 46;
			10409: Pixel = 45;
			10410: Pixel = 62;
			10411: Pixel = 63;
			10412: Pixel = 56;
			10413: Pixel = 41;
			10414: Pixel = 81;
			10415: Pixel = 55;
			10416: Pixel = 22;
			10417: Pixel = 81;
			10418: Pixel = 139;
			10419: Pixel = 121;
			10420: Pixel = 152;
			10421: Pixel = 166;
			10422: Pixel = 159;
			10423: Pixel = 177;
			10424: Pixel = 187;
			10425: Pixel = 188;
			10426: Pixel = 155;
			10427: Pixel = 157;
			10428: Pixel = 188;
			10429: Pixel = 166;
			10430: Pixel = 154;
			10431: Pixel = 157;
			10432: Pixel = 157;
			10433: Pixel = 162;
			10434: Pixel = 168;
			10435: Pixel = 173;
			10436: Pixel = 174;
			10437: Pixel = 177;
			10438: Pixel = 182;
			10439: Pixel = 191;
			10440: Pixel = 195;
			10441: Pixel = 198;
			10442: Pixel = 198;
			10443: Pixel = 200;
			10444: Pixel = 202;
			10445: Pixel = 205;
			10446: Pixel = 208;
			10447: Pixel = 211;
			10448: Pixel = 213;
			10449: Pixel = 208;
			10450: Pixel = 174;
			10451: Pixel = 115;
			10452: Pixel = 80;
			10453: Pixel = 48;
			10454: Pixel = 38;
			10455: Pixel = 56;
			10456: Pixel = 121;
			10457: Pixel = 166;
			10458: Pixel = 74;
			10459: Pixel = 48;
			10460: Pixel = 51;
			10461: Pixel = 57;
			10462: Pixel = 59;
			10463: Pixel = 62;
			10464: Pixel = 63;
			10465: Pixel = 53;
			10466: Pixel = 48;
			10467: Pixel = 50;
			10468: Pixel = 54;
			10469: Pixel = 43;
			10470: Pixel = 55;
			10471: Pixel = 118;
			10472: Pixel = 143;
			10473: Pixel = 134;
			10474: Pixel = 148;
			10475: Pixel = 165;
			10476: Pixel = 162;
			10477: Pixel = 161;
			10478: Pixel = 161;
			10479: Pixel = 159;
			10480: Pixel = 164;
			10481: Pixel = 162;
			10482: Pixel = 161;
			10483: Pixel = 159;
			10484: Pixel = 155;
			10485: Pixel = 154;
			10486: Pixel = 149;
			10487: Pixel = 144;
			10488: Pixel = 147;
			10489: Pixel = 146;
			10490: Pixel = 143;
			10491: Pixel = 144;
			10492: Pixel = 143;
			10493: Pixel = 146;
			10494: Pixel = 149;
			10495: Pixel = 150;
			10496: Pixel = 153;
			10497: Pixel = 153;
			10498: Pixel = 151;
			10499: Pixel = 150;
			10500: Pixel = 102;
			10501: Pixel = 102;
			10502: Pixel = 101;
			10503: Pixel = 99;
			10504: Pixel = 96;
			10505: Pixel = 98;
			10506: Pixel = 91;
			10507: Pixel = 93;
			10508: Pixel = 121;
			10509: Pixel = 147;
			10510: Pixel = 161;
			10511: Pixel = 171;
			10512: Pixel = 173;
			10513: Pixel = 175;
			10514: Pixel = 176;
			10515: Pixel = 174;
			10516: Pixel = 162;
			10517: Pixel = 143;
			10518: Pixel = 110;
			10519: Pixel = 80;
			10520: Pixel = 76;
			10521: Pixel = 85;
			10522: Pixel = 93;
			10523: Pixel = 99;
			10524: Pixel = 101;
			10525: Pixel = 101;
			10526: Pixel = 103;
			10527: Pixel = 104;
			10528: Pixel = 103;
			10529: Pixel = 103;
			10530: Pixel = 104;
			10531: Pixel = 108;
			10532: Pixel = 112;
			10533: Pixel = 117;
			10534: Pixel = 118;
			10535: Pixel = 118;
			10536: Pixel = 117;
			10537: Pixel = 108;
			10538: Pixel = 132;
			10539: Pixel = 118;
			10540: Pixel = 129;
			10541: Pixel = 143;
			10542: Pixel = 118;
			10543: Pixel = 130;
			10544: Pixel = 126;
			10545: Pixel = 124;
			10546: Pixel = 101;
			10547: Pixel = 53;
			10548: Pixel = 84;
			10549: Pixel = 32;
			10550: Pixel = 75;
			10551: Pixel = 79;
			10552: Pixel = 44;
			10553: Pixel = 49;
			10554: Pixel = 61;
			10555: Pixel = 91;
			10556: Pixel = 79;
			10557: Pixel = 41;
			10558: Pixel = 48;
			10559: Pixel = 47;
			10560: Pixel = 71;
			10561: Pixel = 48;
			10562: Pixel = 78;
			10563: Pixel = 50;
			10564: Pixel = 80;
			10565: Pixel = 50;
			10566: Pixel = 31;
			10567: Pixel = 104;
			10568: Pixel = 106;
			10569: Pixel = 144;
			10570: Pixel = 172;
			10571: Pixel = 162;
			10572: Pixel = 159;
			10573: Pixel = 171;
			10574: Pixel = 189;
			10575: Pixel = 185;
			10576: Pixel = 177;
			10577: Pixel = 182;
			10578: Pixel = 172;
			10579: Pixel = 155;
			10580: Pixel = 160;
			10581: Pixel = 166;
			10582: Pixel = 165;
			10583: Pixel = 165;
			10584: Pixel = 171;
			10585: Pixel = 176;
			10586: Pixel = 176;
			10587: Pixel = 177;
			10588: Pixel = 179;
			10589: Pixel = 187;
			10590: Pixel = 194;
			10591: Pixel = 196;
			10592: Pixel = 194;
			10593: Pixel = 197;
			10594: Pixel = 201;
			10595: Pixel = 203;
			10596: Pixel = 206;
			10597: Pixel = 209;
			10598: Pixel = 211;
			10599: Pixel = 208;
			10600: Pixel = 188;
			10601: Pixel = 124;
			10602: Pixel = 83;
			10603: Pixel = 45;
			10604: Pixel = 39;
			10605: Pixel = 51;
			10606: Pixel = 101;
			10607: Pixel = 172;
			10608: Pixel = 88;
			10609: Pixel = 51;
			10610: Pixel = 61;
			10611: Pixel = 60;
			10612: Pixel = 58;
			10613: Pixel = 63;
			10614: Pixel = 63;
			10615: Pixel = 51;
			10616: Pixel = 50;
			10617: Pixel = 52;
			10618: Pixel = 52;
			10619: Pixel = 42;
			10620: Pixel = 75;
			10621: Pixel = 135;
			10622: Pixel = 136;
			10623: Pixel = 133;
			10624: Pixel = 156;
			10625: Pixel = 163;
			10626: Pixel = 162;
			10627: Pixel = 161;
			10628: Pixel = 160;
			10629: Pixel = 160;
			10630: Pixel = 162;
			10631: Pixel = 164;
			10632: Pixel = 166;
			10633: Pixel = 165;
			10634: Pixel = 159;
			10635: Pixel = 156;
			10636: Pixel = 153;
			10637: Pixel = 148;
			10638: Pixel = 147;
			10639: Pixel = 146;
			10640: Pixel = 144;
			10641: Pixel = 143;
			10642: Pixel = 142;
			10643: Pixel = 142;
			10644: Pixel = 142;
			10645: Pixel = 143;
			10646: Pixel = 148;
			10647: Pixel = 148;
			10648: Pixel = 150;
			10649: Pixel = 152;
			10650: Pixel = 101;
			10651: Pixel = 101;
			10652: Pixel = 98;
			10653: Pixel = 98;
			10654: Pixel = 98;
			10655: Pixel = 97;
			10656: Pixel = 92;
			10657: Pixel = 93;
			10658: Pixel = 120;
			10659: Pixel = 145;
			10660: Pixel = 160;
			10661: Pixel = 169;
			10662: Pixel = 173;
			10663: Pixel = 175;
			10664: Pixel = 176;
			10665: Pixel = 174;
			10666: Pixel = 162;
			10667: Pixel = 144;
			10668: Pixel = 111;
			10669: Pixel = 79;
			10670: Pixel = 77;
			10671: Pixel = 86;
			10672: Pixel = 92;
			10673: Pixel = 98;
			10674: Pixel = 102;
			10675: Pixel = 102;
			10676: Pixel = 102;
			10677: Pixel = 101;
			10678: Pixel = 101;
			10679: Pixel = 101;
			10680: Pixel = 104;
			10681: Pixel = 109;
			10682: Pixel = 113;
			10683: Pixel = 115;
			10684: Pixel = 118;
			10685: Pixel = 120;
			10686: Pixel = 120;
			10687: Pixel = 148;
			10688: Pixel = 151;
			10689: Pixel = 95;
			10690: Pixel = 91;
			10691: Pixel = 126;
			10692: Pixel = 125;
			10693: Pixel = 128;
			10694: Pixel = 122;
			10695: Pixel = 118;
			10696: Pixel = 66;
			10697: Pixel = 72;
			10698: Pixel = 80;
			10699: Pixel = 28;
			10700: Pixel = 91;
			10701: Pixel = 72;
			10702: Pixel = 36;
			10703: Pixel = 54;
			10704: Pixel = 73;
			10705: Pixel = 70;
			10706: Pixel = 48;
			10707: Pixel = 41;
			10708: Pixel = 49;
			10709: Pixel = 55;
			10710: Pixel = 57;
			10711: Pixel = 48;
			10712: Pixel = 83;
			10713: Pixel = 58;
			10714: Pixel = 70;
			10715: Pixel = 34;
			10716: Pixel = 93;
			10717: Pixel = 126;
			10718: Pixel = 127;
			10719: Pixel = 180;
			10720: Pixel = 170;
			10721: Pixel = 176;
			10722: Pixel = 155;
			10723: Pixel = 171;
			10724: Pixel = 191;
			10725: Pixel = 190;
			10726: Pixel = 189;
			10727: Pixel = 145;
			10728: Pixel = 98;
			10729: Pixel = 116;
			10730: Pixel = 136;
			10731: Pixel = 149;
			10732: Pixel = 160;
			10733: Pixel = 172;
			10734: Pixel = 177;
			10735: Pixel = 178;
			10736: Pixel = 179;
			10737: Pixel = 175;
			10738: Pixel = 178;
			10739: Pixel = 182;
			10740: Pixel = 190;
			10741: Pixel = 196;
			10742: Pixel = 193;
			10743: Pixel = 194;
			10744: Pixel = 197;
			10745: Pixel = 201;
			10746: Pixel = 202;
			10747: Pixel = 206;
			10748: Pixel = 210;
			10749: Pixel = 207;
			10750: Pixel = 186;
			10751: Pixel = 123;
			10752: Pixel = 62;
			10753: Pixel = 44;
			10754: Pixel = 39;
			10755: Pixel = 47;
			10756: Pixel = 86;
			10757: Pixel = 174;
			10758: Pixel = 101;
			10759: Pixel = 57;
			10760: Pixel = 64;
			10761: Pixel = 60;
			10762: Pixel = 61;
			10763: Pixel = 69;
			10764: Pixel = 59;
			10765: Pixel = 48;
			10766: Pixel = 51;
			10767: Pixel = 54;
			10768: Pixel = 50;
			10769: Pixel = 48;
			10770: Pixel = 101;
			10771: Pixel = 140;
			10772: Pixel = 132;
			10773: Pixel = 139;
			10774: Pixel = 160;
			10775: Pixel = 160;
			10776: Pixel = 160;
			10777: Pixel = 160;
			10778: Pixel = 160;
			10779: Pixel = 159;
			10780: Pixel = 159;
			10781: Pixel = 162;
			10782: Pixel = 163;
			10783: Pixel = 164;
			10784: Pixel = 161;
			10785: Pixel = 157;
			10786: Pixel = 156;
			10787: Pixel = 154;
			10788: Pixel = 151;
			10789: Pixel = 149;
			10790: Pixel = 146;
			10791: Pixel = 145;
			10792: Pixel = 146;
			10793: Pixel = 144;
			10794: Pixel = 142;
			10795: Pixel = 140;
			10796: Pixel = 142;
			10797: Pixel = 141;
			10798: Pixel = 142;
			10799: Pixel = 144;
			10800: Pixel = 100;
			10801: Pixel = 100;
			10802: Pixel = 100;
			10803: Pixel = 100;
			10804: Pixel = 100;
			10805: Pixel = 99;
			10806: Pixel = 93;
			10807: Pixel = 92;
			10808: Pixel = 120;
			10809: Pixel = 145;
			10810: Pixel = 161;
			10811: Pixel = 170;
			10812: Pixel = 175;
			10813: Pixel = 176;
			10814: Pixel = 176;
			10815: Pixel = 173;
			10816: Pixel = 163;
			10817: Pixel = 145;
			10818: Pixel = 111;
			10819: Pixel = 79;
			10820: Pixel = 77;
			10821: Pixel = 86;
			10822: Pixel = 92;
			10823: Pixel = 96;
			10824: Pixel = 102;
			10825: Pixel = 103;
			10826: Pixel = 101;
			10827: Pixel = 103;
			10828: Pixel = 102;
			10829: Pixel = 101;
			10830: Pixel = 104;
			10831: Pixel = 107;
			10832: Pixel = 115;
			10833: Pixel = 118;
			10834: Pixel = 119;
			10835: Pixel = 117;
			10836: Pixel = 131;
			10837: Pixel = 188;
			10838: Pixel = 92;
			10839: Pixel = 38;
			10840: Pixel = 30;
			10841: Pixel = 94;
			10842: Pixel = 182;
			10843: Pixel = 138;
			10844: Pixel = 91;
			10845: Pixel = 76;
			10846: Pixel = 55;
			10847: Pixel = 101;
			10848: Pixel = 54;
			10849: Pixel = 42;
			10850: Pixel = 119;
			10851: Pixel = 58;
			10852: Pixel = 38;
			10853: Pixel = 52;
			10854: Pixel = 56;
			10855: Pixel = 54;
			10856: Pixel = 49;
			10857: Pixel = 49;
			10858: Pixel = 46;
			10859: Pixel = 57;
			10860: Pixel = 71;
			10861: Pixel = 58;
			10862: Pixel = 76;
			10863: Pixel = 63;
			10864: Pixel = 39;
			10865: Pixel = 60;
			10866: Pixel = 132;
			10867: Pixel = 113;
			10868: Pixel = 177;
			10869: Pixel = 171;
			10870: Pixel = 188;
			10871: Pixel = 176;
			10872: Pixel = 151;
			10873: Pixel = 176;
			10874: Pixel = 196;
			10875: Pixel = 195;
			10876: Pixel = 145;
			10877: Pixel = 105;
			10878: Pixel = 114;
			10879: Pixel = 109;
			10880: Pixel = 98;
			10881: Pixel = 83;
			10882: Pixel = 94;
			10883: Pixel = 122;
			10884: Pixel = 157;
			10885: Pixel = 181;
			10886: Pixel = 179;
			10887: Pixel = 176;
			10888: Pixel = 174;
			10889: Pixel = 176;
			10890: Pixel = 187;
			10891: Pixel = 194;
			10892: Pixel = 190;
			10893: Pixel = 189;
			10894: Pixel = 193;
			10895: Pixel = 198;
			10896: Pixel = 202;
			10897: Pixel = 209;
			10898: Pixel = 200;
			10899: Pixel = 169;
			10900: Pixel = 131;
			10901: Pixel = 85;
			10902: Pixel = 52;
			10903: Pixel = 42;
			10904: Pixel = 37;
			10905: Pixel = 50;
			10906: Pixel = 71;
			10907: Pixel = 168;
			10908: Pixel = 122;
			10909: Pixel = 49;
			10910: Pixel = 64;
			10911: Pixel = 60;
			10912: Pixel = 62;
			10913: Pixel = 65;
			10914: Pixel = 54;
			10915: Pixel = 48;
			10916: Pixel = 50;
			10917: Pixel = 54;
			10918: Pixel = 46;
			10919: Pixel = 57;
			10920: Pixel = 119;
			10921: Pixel = 141;
			10922: Pixel = 129;
			10923: Pixel = 148;
			10924: Pixel = 163;
			10925: Pixel = 159;
			10926: Pixel = 158;
			10927: Pixel = 157;
			10928: Pixel = 158;
			10929: Pixel = 157;
			10930: Pixel = 157;
			10931: Pixel = 157;
			10932: Pixel = 159;
			10933: Pixel = 159;
			10934: Pixel = 161;
			10935: Pixel = 157;
			10936: Pixel = 153;
			10937: Pixel = 156;
			10938: Pixel = 155;
			10939: Pixel = 153;
			10940: Pixel = 152;
			10941: Pixel = 152;
			10942: Pixel = 151;
			10943: Pixel = 148;
			10944: Pixel = 142;
			10945: Pixel = 141;
			10946: Pixel = 141;
			10947: Pixel = 140;
			10948: Pixel = 136;
			10949: Pixel = 134;
			10950: Pixel = 103;
			10951: Pixel = 102;
			10952: Pixel = 102;
			10953: Pixel = 101;
			10954: Pixel = 100;
			10955: Pixel = 99;
			10956: Pixel = 93;
			10957: Pixel = 91;
			10958: Pixel = 118;
			10959: Pixel = 145;
			10960: Pixel = 159;
			10961: Pixel = 172;
			10962: Pixel = 174;
			10963: Pixel = 175;
			10964: Pixel = 177;
			10965: Pixel = 175;
			10966: Pixel = 163;
			10967: Pixel = 146;
			10968: Pixel = 112;
			10969: Pixel = 78;
			10970: Pixel = 80;
			10971: Pixel = 86;
			10972: Pixel = 93;
			10973: Pixel = 96;
			10974: Pixel = 103;
			10975: Pixel = 103;
			10976: Pixel = 101;
			10977: Pixel = 99;
			10978: Pixel = 100;
			10979: Pixel = 101;
			10980: Pixel = 102;
			10981: Pixel = 107;
			10982: Pixel = 112;
			10983: Pixel = 114;
			10984: Pixel = 117;
			10985: Pixel = 131;
			10986: Pixel = 138;
			10987: Pixel = 153;
			10988: Pixel = 88;
			10989: Pixel = 40;
			10990: Pixel = 36;
			10991: Pixel = 120;
			10992: Pixel = 134;
			10993: Pixel = 96;
			10994: Pixel = 77;
			10995: Pixel = 64;
			10996: Pixel = 78;
			10997: Pixel = 79;
			10998: Pixel = 42;
			10999: Pixel = 78;
			11000: Pixel = 100;
			11001: Pixel = 70;
			11002: Pixel = 32;
			11003: Pixel = 65;
			11004: Pixel = 63;
			11005: Pixel = 64;
			11006: Pixel = 71;
			11007: Pixel = 48;
			11008: Pixel = 40;
			11009: Pixel = 37;
			11010: Pixel = 72;
			11011: Pixel = 90;
			11012: Pixel = 66;
			11013: Pixel = 54;
			11014: Pixel = 33;
			11015: Pixel = 132;
			11016: Pixel = 123;
			11017: Pixel = 166;
			11018: Pixel = 171;
			11019: Pixel = 183;
			11020: Pixel = 195;
			11021: Pixel = 159;
			11022: Pixel = 161;
			11023: Pixel = 195;
			11024: Pixel = 189;
			11025: Pixel = 136;
			11026: Pixel = 129;
			11027: Pixel = 155;
			11028: Pixel = 151;
			11029: Pixel = 157;
			11030: Pixel = 142;
			11031: Pixel = 107;
			11032: Pixel = 76;
			11033: Pixel = 67;
			11034: Pixel = 77;
			11035: Pixel = 122;
			11036: Pixel = 165;
			11037: Pixel = 172;
			11038: Pixel = 170;
			11039: Pixel = 174;
			11040: Pixel = 184;
			11041: Pixel = 192;
			11042: Pixel = 189;
			11043: Pixel = 189;
			11044: Pixel = 191;
			11045: Pixel = 192;
			11046: Pixel = 182;
			11047: Pixel = 146;
			11048: Pixel = 114;
			11049: Pixel = 93;
			11050: Pixel = 96;
			11051: Pixel = 101;
			11052: Pixel = 86;
			11053: Pixel = 53;
			11054: Pixel = 42;
			11055: Pixel = 46;
			11056: Pixel = 61;
			11057: Pixel = 161;
			11058: Pixel = 137;
			11059: Pixel = 56;
			11060: Pixel = 59;
			11061: Pixel = 68;
			11062: Pixel = 65;
			11063: Pixel = 60;
			11064: Pixel = 50;
			11065: Pixel = 49;
			11066: Pixel = 49;
			11067: Pixel = 58;
			11068: Pixel = 49;
			11069: Pixel = 70;
			11070: Pixel = 135;
			11071: Pixel = 134;
			11072: Pixel = 132;
			11073: Pixel = 157;
			11074: Pixel = 163;
			11075: Pixel = 159;
			11076: Pixel = 158;
			11077: Pixel = 157;
			11078: Pixel = 157;
			11079: Pixel = 156;
			11080: Pixel = 155;
			11081: Pixel = 155;
			11082: Pixel = 156;
			11083: Pixel = 158;
			11084: Pixel = 158;
			11085: Pixel = 155;
			11086: Pixel = 154;
			11087: Pixel = 154;
			11088: Pixel = 154;
			11089: Pixel = 154;
			11090: Pixel = 155;
			11091: Pixel = 156;
			11092: Pixel = 154;
			11093: Pixel = 152;
			11094: Pixel = 148;
			11095: Pixel = 144;
			11096: Pixel = 142;
			11097: Pixel = 139;
			11098: Pixel = 134;
			11099: Pixel = 132;
			11100: Pixel = 99;
			11101: Pixel = 101;
			11102: Pixel = 104;
			11103: Pixel = 104;
			11104: Pixel = 100;
			11105: Pixel = 98;
			11106: Pixel = 89;
			11107: Pixel = 90;
			11108: Pixel = 118;
			11109: Pixel = 144;
			11110: Pixel = 158;
			11111: Pixel = 172;
			11112: Pixel = 174;
			11113: Pixel = 174;
			11114: Pixel = 176;
			11115: Pixel = 177;
			11116: Pixel = 164;
			11117: Pixel = 147;
			11118: Pixel = 114;
			11119: Pixel = 79;
			11120: Pixel = 79;
			11121: Pixel = 87;
			11122: Pixel = 94;
			11123: Pixel = 99;
			11124: Pixel = 103;
			11125: Pixel = 101;
			11126: Pixel = 101;
			11127: Pixel = 100;
			11128: Pixel = 98;
			11129: Pixel = 100;
			11130: Pixel = 101;
			11131: Pixel = 105;
			11132: Pixel = 105;
			11133: Pixel = 106;
			11134: Pixel = 127;
			11135: Pixel = 157;
			11136: Pixel = 148;
			11137: Pixel = 152;
			11138: Pixel = 138;
			11139: Pixel = 117;
			11140: Pixel = 93;
			11141: Pixel = 114;
			11142: Pixel = 122;
			11143: Pixel = 72;
			11144: Pixel = 59;
			11145: Pixel = 61;
			11146: Pixel = 102;
			11147: Pixel = 62;
			11148: Pixel = 78;
			11149: Pixel = 81;
			11150: Pixel = 51;
			11151: Pixel = 92;
			11152: Pixel = 39;
			11153: Pixel = 69;
			11154: Pixel = 44;
			11155: Pixel = 47;
			11156: Pixel = 97;
			11157: Pixel = 47;
			11158: Pixel = 37;
			11159: Pixel = 45;
			11160: Pixel = 41;
			11161: Pixel = 69;
			11162: Pixel = 65;
			11163: Pixel = 27;
			11164: Pixel = 91;
			11165: Pixel = 132;
			11166: Pixel = 157;
			11167: Pixel = 176;
			11168: Pixel = 175;
			11169: Pixel = 197;
			11170: Pixel = 185;
			11171: Pixel = 157;
			11172: Pixel = 192;
			11173: Pixel = 182;
			11174: Pixel = 115;
			11175: Pixel = 111;
			11176: Pixel = 118;
			11177: Pixel = 126;
			11178: Pixel = 94;
			11179: Pixel = 123;
			11180: Pixel = 136;
			11181: Pixel = 109;
			11182: Pixel = 113;
			11183: Pixel = 104;
			11184: Pixel = 92;
			11185: Pixel = 93;
			11186: Pixel = 132;
			11187: Pixel = 159;
			11188: Pixel = 162;
			11189: Pixel = 167;
			11190: Pixel = 181;
			11191: Pixel = 192;
			11192: Pixel = 193;
			11193: Pixel = 189;
			11194: Pixel = 186;
			11195: Pixel = 172;
			11196: Pixel = 132;
			11197: Pixel = 101;
			11198: Pixel = 102;
			11199: Pixel = 96;
			11200: Pixel = 110;
			11201: Pixel = 104;
			11202: Pixel = 85;
			11203: Pixel = 66;
			11204: Pixel = 47;
			11205: Pixel = 45;
			11206: Pixel = 61;
			11207: Pixel = 153;
			11208: Pixel = 140;
			11209: Pixel = 64;
			11210: Pixel = 52;
			11211: Pixel = 65;
			11212: Pixel = 63;
			11213: Pixel = 60;
			11214: Pixel = 48;
			11215: Pixel = 51;
			11216: Pixel = 53;
			11217: Pixel = 53;
			11218: Pixel = 52;
			11219: Pixel = 93;
			11220: Pixel = 140;
			11221: Pixel = 128;
			11222: Pixel = 140;
			11223: Pixel = 160;
			11224: Pixel = 160;
			11225: Pixel = 158;
			11226: Pixel = 157;
			11227: Pixel = 156;
			11228: Pixel = 157;
			11229: Pixel = 155;
			11230: Pixel = 154;
			11231: Pixel = 154;
			11232: Pixel = 156;
			11233: Pixel = 158;
			11234: Pixel = 157;
			11235: Pixel = 155;
			11236: Pixel = 155;
			11237: Pixel = 153;
			11238: Pixel = 153;
			11239: Pixel = 154;
			11240: Pixel = 154;
			11241: Pixel = 156;
			11242: Pixel = 156;
			11243: Pixel = 154;
			11244: Pixel = 150;
			11245: Pixel = 151;
			11246: Pixel = 147;
			11247: Pixel = 140;
			11248: Pixel = 136;
			11249: Pixel = 132;
			11250: Pixel = 101;
			11251: Pixel = 102;
			11252: Pixel = 102;
			11253: Pixel = 100;
			11254: Pixel = 99;
			11255: Pixel = 96;
			11256: Pixel = 87;
			11257: Pixel = 88;
			11258: Pixel = 120;
			11259: Pixel = 144;
			11260: Pixel = 159;
			11261: Pixel = 171;
			11262: Pixel = 176;
			11263: Pixel = 176;
			11264: Pixel = 177;
			11265: Pixel = 174;
			11266: Pixel = 164;
			11267: Pixel = 149;
			11268: Pixel = 115;
			11269: Pixel = 80;
			11270: Pixel = 76;
			11271: Pixel = 84;
			11272: Pixel = 91;
			11273: Pixel = 98;
			11274: Pixel = 101;
			11275: Pixel = 102;
			11276: Pixel = 100;
			11277: Pixel = 99;
			11278: Pixel = 99;
			11279: Pixel = 98;
			11280: Pixel = 98;
			11281: Pixel = 96;
			11282: Pixel = 119;
			11283: Pixel = 142;
			11284: Pixel = 143;
			11285: Pixel = 153;
			11286: Pixel = 153;
			11287: Pixel = 157;
			11288: Pixel = 159;
			11289: Pixel = 154;
			11290: Pixel = 134;
			11291: Pixel = 63;
			11292: Pixel = 49;
			11293: Pixel = 61;
			11294: Pixel = 67;
			11295: Pixel = 105;
			11296: Pixel = 88;
			11297: Pixel = 68;
			11298: Pixel = 99;
			11299: Pixel = 66;
			11300: Pixel = 38;
			11301: Pixel = 81;
			11302: Pixel = 48;
			11303: Pixel = 71;
			11304: Pixel = 45;
			11305: Pixel = 34;
			11306: Pixel = 80;
			11307: Pixel = 88;
			11308: Pixel = 38;
			11309: Pixel = 42;
			11310: Pixel = 46;
			11311: Pixel = 37;
			11312: Pixel = 37;
			11313: Pixel = 54;
			11314: Pixel = 134;
			11315: Pixel = 134;
			11316: Pixel = 181;
			11317: Pixel = 170;
			11318: Pixel = 192;
			11319: Pixel = 201;
			11320: Pixel = 180;
			11321: Pixel = 189;
			11322: Pixel = 170;
			11323: Pixel = 86;
			11324: Pixel = 77;
			11325: Pixel = 77;
			11326: Pixel = 65;
			11327: Pixel = 60;
			11328: Pixel = 49;
			11329: Pixel = 55;
			11330: Pixel = 51;
			11331: Pixel = 45;
			11332: Pixel = 77;
			11333: Pixel = 119;
			11334: Pixel = 132;
			11335: Pixel = 122;
			11336: Pixel = 127;
			11337: Pixel = 145;
			11338: Pixel = 155;
			11339: Pixel = 160;
			11340: Pixel = 181;
			11341: Pixel = 195;
			11342: Pixel = 196;
			11343: Pixel = 194;
			11344: Pixel = 188;
			11345: Pixel = 137;
			11346: Pixel = 98;
			11347: Pixel = 77;
			11348: Pixel = 58;
			11349: Pixel = 49;
			11350: Pixel = 57;
			11351: Pixel = 59;
			11352: Pixel = 66;
			11353: Pixel = 63;
			11354: Pixel = 42;
			11355: Pixel = 44;
			11356: Pixel = 62;
			11357: Pixel = 148;
			11358: Pixel = 143;
			11359: Pixel = 78;
			11360: Pixel = 53;
			11361: Pixel = 68;
			11362: Pixel = 62;
			11363: Pixel = 52;
			11364: Pixel = 48;
			11365: Pixel = 49;
			11366: Pixel = 53;
			11367: Pixel = 47;
			11368: Pixel = 47;
			11369: Pixel = 118;
			11370: Pixel = 141;
			11371: Pixel = 129;
			11372: Pixel = 148;
			11373: Pixel = 161;
			11374: Pixel = 158;
			11375: Pixel = 157;
			11376: Pixel = 155;
			11377: Pixel = 155;
			11378: Pixel = 156;
			11379: Pixel = 156;
			11380: Pixel = 154;
			11381: Pixel = 155;
			11382: Pixel = 155;
			11383: Pixel = 156;
			11384: Pixel = 157;
			11385: Pixel = 154;
			11386: Pixel = 153;
			11387: Pixel = 152;
			11388: Pixel = 154;
			11389: Pixel = 152;
			11390: Pixel = 153;
			11391: Pixel = 154;
			11392: Pixel = 155;
			11393: Pixel = 152;
			11394: Pixel = 147;
			11395: Pixel = 147;
			11396: Pixel = 146;
			11397: Pixel = 143;
			11398: Pixel = 139;
			11399: Pixel = 135;
			11400: Pixel = 97;
			11401: Pixel = 97;
			11402: Pixel = 96;
			11403: Pixel = 96;
			11404: Pixel = 94;
			11405: Pixel = 93;
			11406: Pixel = 83;
			11407: Pixel = 82;
			11408: Pixel = 113;
			11409: Pixel = 142;
			11410: Pixel = 159;
			11411: Pixel = 171;
			11412: Pixel = 175;
			11413: Pixel = 177;
			11414: Pixel = 177;
			11415: Pixel = 174;
			11416: Pixel = 161;
			11417: Pixel = 146;
			11418: Pixel = 114;
			11419: Pixel = 79;
			11420: Pixel = 73;
			11421: Pixel = 84;
			11422: Pixel = 88;
			11423: Pixel = 93;
			11424: Pixel = 99;
			11425: Pixel = 101;
			11426: Pixel = 98;
			11427: Pixel = 97;
			11428: Pixel = 97;
			11429: Pixel = 95;
			11430: Pixel = 86;
			11431: Pixel = 123;
			11432: Pixel = 185;
			11433: Pixel = 170;
			11434: Pixel = 137;
			11435: Pixel = 150;
			11436: Pixel = 153;
			11437: Pixel = 150;
			11438: Pixel = 117;
			11439: Pixel = 70;
			11440: Pixel = 74;
			11441: Pixel = 26;
			11442: Pixel = 57;
			11443: Pixel = 98;
			11444: Pixel = 82;
			11445: Pixel = 101;
			11446: Pixel = 79;
			11447: Pixel = 78;
			11448: Pixel = 112;
			11449: Pixel = 70;
			11450: Pixel = 44;
			11451: Pixel = 64;
			11452: Pixel = 58;
			11453: Pixel = 83;
			11454: Pixel = 50;
			11455: Pixel = 37;
			11456: Pixel = 38;
			11457: Pixel = 98;
			11458: Pixel = 98;
			11459: Pixel = 48;
			11460: Pixel = 43;
			11461: Pixel = 40;
			11462: Pixel = 28;
			11463: Pixel = 114;
			11464: Pixel = 131;
			11465: Pixel = 175;
			11466: Pixel = 171;
			11467: Pixel = 179;
			11468: Pixel = 198;
			11469: Pixel = 192;
			11470: Pixel = 195;
			11471: Pixel = 169;
			11472: Pixel = 75;
			11473: Pixel = 59;
			11474: Pixel = 52;
			11475: Pixel = 47;
			11476: Pixel = 49;
			11477: Pixel = 45;
			11478: Pixel = 45;
			11479: Pixel = 76;
			11480: Pixel = 94;
			11481: Pixel = 45;
			11482: Pixel = 31;
			11483: Pixel = 65;
			11484: Pixel = 128;
			11485: Pixel = 132;
			11486: Pixel = 130;
			11487: Pixel = 140;
			11488: Pixel = 149;
			11489: Pixel = 160;
			11490: Pixel = 181;
			11491: Pixel = 198;
			11492: Pixel = 204;
			11493: Pixel = 201;
			11494: Pixel = 124;
			11495: Pixel = 62;
			11496: Pixel = 49;
			11497: Pixel = 53;
			11498: Pixel = 75;
			11499: Pixel = 53;
			11500: Pixel = 48;
			11501: Pixel = 57;
			11502: Pixel = 58;
			11503: Pixel = 51;
			11504: Pixel = 43;
			11505: Pixel = 45;
			11506: Pixel = 57;
			11507: Pixel = 143;
			11508: Pixel = 146;
			11509: Pixel = 78;
			11510: Pixel = 60;
			11511: Pixel = 67;
			11512: Pixel = 59;
			11513: Pixel = 48;
			11514: Pixel = 48;
			11515: Pixel = 50;
			11516: Pixel = 56;
			11517: Pixel = 45;
			11518: Pixel = 57;
			11519: Pixel = 133;
			11520: Pixel = 138;
			11521: Pixel = 137;
			11522: Pixel = 158;
			11523: Pixel = 159;
			11524: Pixel = 156;
			11525: Pixel = 155;
			11526: Pixel = 153;
			11527: Pixel = 153;
			11528: Pixel = 153;
			11529: Pixel = 153;
			11530: Pixel = 156;
			11531: Pixel = 155;
			11532: Pixel = 154;
			11533: Pixel = 156;
			11534: Pixel = 155;
			11535: Pixel = 154;
			11536: Pixel = 152;
			11537: Pixel = 154;
			11538: Pixel = 153;
			11539: Pixel = 152;
			11540: Pixel = 151;
			11541: Pixel = 152;
			11542: Pixel = 151;
			11543: Pixel = 147;
			11544: Pixel = 145;
			11545: Pixel = 142;
			11546: Pixel = 141;
			11547: Pixel = 140;
			11548: Pixel = 139;
			11549: Pixel = 136;
			11550: Pixel = 96;
			11551: Pixel = 96;
			11552: Pixel = 93;
			11553: Pixel = 93;
			11554: Pixel = 91;
			11555: Pixel = 87;
			11556: Pixel = 79;
			11557: Pixel = 77;
			11558: Pixel = 112;
			11559: Pixel = 142;
			11560: Pixel = 159;
			11561: Pixel = 174;
			11562: Pixel = 175;
			11563: Pixel = 176;
			11564: Pixel = 177;
			11565: Pixel = 175;
			11566: Pixel = 162;
			11567: Pixel = 144;
			11568: Pixel = 114;
			11569: Pixel = 77;
			11570: Pixel = 74;
			11571: Pixel = 86;
			11572: Pixel = 92;
			11573: Pixel = 96;
			11574: Pixel = 97;
			11575: Pixel = 97;
			11576: Pixel = 97;
			11577: Pixel = 97;
			11578: Pixel = 93;
			11579: Pixel = 89;
			11580: Pixel = 83;
			11581: Pixel = 168;
			11582: Pixel = 207;
			11583: Pixel = 141;
			11584: Pixel = 134;
			11585: Pixel = 153;
			11586: Pixel = 143;
			11587: Pixel = 130;
			11588: Pixel = 111;
			11589: Pixel = 60;
			11590: Pixel = 37;
			11591: Pixel = 56;
			11592: Pixel = 100;
			11593: Pixel = 60;
			11594: Pixel = 82;
			11595: Pixel = 42;
			11596: Pixel = 73;
			11597: Pixel = 101;
			11598: Pixel = 108;
			11599: Pixel = 56;
			11600: Pixel = 45;
			11601: Pixel = 51;
			11602: Pixel = 43;
			11603: Pixel = 87;
			11604: Pixel = 66;
			11605: Pixel = 41;
			11606: Pixel = 41;
			11607: Pixel = 49;
			11608: Pixel = 67;
			11609: Pixel = 72;
			11610: Pixel = 56;
			11611: Pixel = 32;
			11612: Pixel = 74;
			11613: Pixel = 131;
			11614: Pixel = 152;
			11615: Pixel = 183;
			11616: Pixel = 174;
			11617: Pixel = 185;
			11618: Pixel = 199;
			11619: Pixel = 202;
			11620: Pixel = 175;
			11621: Pixel = 85;
			11622: Pixel = 67;
			11623: Pixel = 49;
			11624: Pixel = 50;
			11625: Pixel = 63;
			11626: Pixel = 59;
			11627: Pixel = 46;
			11628: Pixel = 58;
			11629: Pixel = 114;
			11630: Pixel = 200;
			11631: Pixel = 139;
			11632: Pixel = 57;
			11633: Pixel = 62;
			11634: Pixel = 102;
			11635: Pixel = 127;
			11636: Pixel = 125;
			11637: Pixel = 138;
			11638: Pixel = 144;
			11639: Pixel = 157;
			11640: Pixel = 180;
			11641: Pixel = 207;
			11642: Pixel = 218;
			11643: Pixel = 140;
			11644: Pixel = 45;
			11645: Pixel = 43;
			11646: Pixel = 52;
			11647: Pixel = 100;
			11648: Pixel = 148;
			11649: Pixel = 106;
			11650: Pixel = 42;
			11651: Pixel = 51;
			11652: Pixel = 55;
			11653: Pixel = 48;
			11654: Pixel = 45;
			11655: Pixel = 48;
			11656: Pixel = 55;
			11657: Pixel = 138;
			11658: Pixel = 148;
			11659: Pixel = 80;
			11660: Pixel = 67;
			11661: Pixel = 71;
			11662: Pixel = 57;
			11663: Pixel = 47;
			11664: Pixel = 48;
			11665: Pixel = 52;
			11666: Pixel = 49;
			11667: Pixel = 45;
			11668: Pixel = 88;
			11669: Pixel = 144;
			11670: Pixel = 138;
			11671: Pixel = 145;
			11672: Pixel = 160;
			11673: Pixel = 157;
			11674: Pixel = 156;
			11675: Pixel = 155;
			11676: Pixel = 153;
			11677: Pixel = 153;
			11678: Pixel = 153;
			11679: Pixel = 153;
			11680: Pixel = 153;
			11681: Pixel = 153;
			11682: Pixel = 153;
			11683: Pixel = 153;
			11684: Pixel = 153;
			11685: Pixel = 153;
			11686: Pixel = 152;
			11687: Pixel = 153;
			11688: Pixel = 152;
			11689: Pixel = 149;
			11690: Pixel = 148;
			11691: Pixel = 151;
			11692: Pixel = 146;
			11693: Pixel = 143;
			11694: Pixel = 141;
			11695: Pixel = 138;
			11696: Pixel = 135;
			11697: Pixel = 136;
			11698: Pixel = 133;
			11699: Pixel = 131;
			11700: Pixel = 99;
			11701: Pixel = 98;
			11702: Pixel = 96;
			11703: Pixel = 96;
			11704: Pixel = 91;
			11705: Pixel = 86;
			11706: Pixel = 78;
			11707: Pixel = 76;
			11708: Pixel = 113;
			11709: Pixel = 142;
			11710: Pixel = 161;
			11711: Pixel = 174;
			11712: Pixel = 176;
			11713: Pixel = 177;
			11714: Pixel = 180;
			11715: Pixel = 178;
			11716: Pixel = 164;
			11717: Pixel = 143;
			11718: Pixel = 115;
			11719: Pixel = 79;
			11720: Pixel = 77;
			11721: Pixel = 88;
			11722: Pixel = 96;
			11723: Pixel = 100;
			11724: Pixel = 101;
			11725: Pixel = 99;
			11726: Pixel = 101;
			11727: Pixel = 101;
			11728: Pixel = 101;
			11729: Pixel = 97;
			11730: Pixel = 62;
			11731: Pixel = 126;
			11732: Pixel = 142;
			11733: Pixel = 160;
			11734: Pixel = 158;
			11735: Pixel = 155;
			11736: Pixel = 128;
			11737: Pixel = 110;
			11738: Pixel = 69;
			11739: Pixel = 35;
			11740: Pixel = 62;
			11741: Pixel = 92;
			11742: Pixel = 48;
			11743: Pixel = 64;
			11744: Pixel = 68;
			11745: Pixel = 42;
			11746: Pixel = 84;
			11747: Pixel = 105;
			11748: Pixel = 105;
			11749: Pixel = 52;
			11750: Pixel = 45;
			11751: Pixel = 46;
			11752: Pixel = 37;
			11753: Pixel = 66;
			11754: Pixel = 91;
			11755: Pixel = 40;
			11756: Pixel = 43;
			11757: Pixel = 50;
			11758: Pixel = 40;
			11759: Pixel = 43;
			11760: Pixel = 41;
			11761: Pixel = 50;
			11762: Pixel = 110;
			11763: Pixel = 125;
			11764: Pixel = 176;
			11765: Pixel = 161;
			11766: Pixel = 182;
			11767: Pixel = 196;
			11768: Pixel = 204;
			11769: Pixel = 188;
			11770: Pixel = 110;
			11771: Pixel = 98;
			11772: Pixel = 77;
			11773: Pixel = 49;
			11774: Pixel = 59;
			11775: Pixel = 103;
			11776: Pixel = 77;
			11777: Pixel = 73;
			11778: Pixel = 62;
			11779: Pixel = 116;
			11780: Pixel = 212;
			11781: Pixel = 209;
			11782: Pixel = 130;
			11783: Pixel = 95;
			11784: Pixel = 106;
			11785: Pixel = 110;
			11786: Pixel = 119;
			11787: Pixel = 131;
			11788: Pixel = 141;
			11789: Pixel = 159;
			11790: Pixel = 186;
			11791: Pixel = 218;
			11792: Pixel = 193;
			11793: Pixel = 95;
			11794: Pixel = 71;
			11795: Pixel = 74;
			11796: Pixel = 71;
			11797: Pixel = 76;
			11798: Pixel = 156;
			11799: Pixel = 137;
			11800: Pixel = 58;
			11801: Pixel = 44;
			11802: Pixel = 46;
			11803: Pixel = 47;
			11804: Pixel = 45;
			11805: Pixel = 55;
			11806: Pixel = 57;
			11807: Pixel = 132;
			11808: Pixel = 156;
			11809: Pixel = 84;
			11810: Pixel = 79;
			11811: Pixel = 67;
			11812: Pixel = 53;
			11813: Pixel = 48;
			11814: Pixel = 51;
			11815: Pixel = 52;
			11816: Pixel = 46;
			11817: Pixel = 53;
			11818: Pixel = 113;
			11819: Pixel = 144;
			11820: Pixel = 135;
			11821: Pixel = 150;
			11822: Pixel = 159;
			11823: Pixel = 156;
			11824: Pixel = 157;
			11825: Pixel = 155;
			11826: Pixel = 151;
			11827: Pixel = 152;
			11828: Pixel = 152;
			11829: Pixel = 151;
			11830: Pixel = 152;
			11831: Pixel = 153;
			11832: Pixel = 152;
			11833: Pixel = 151;
			11834: Pixel = 153;
			11835: Pixel = 152;
			11836: Pixel = 151;
			11837: Pixel = 149;
			11838: Pixel = 149;
			11839: Pixel = 147;
			11840: Pixel = 146;
			11841: Pixel = 146;
			11842: Pixel = 142;
			11843: Pixel = 141;
			11844: Pixel = 138;
			11845: Pixel = 132;
			11846: Pixel = 129;
			11847: Pixel = 128;
			11848: Pixel = 131;
			11849: Pixel = 141;
			11850: Pixel = 99;
			11851: Pixel = 98;
			11852: Pixel = 97;
			11853: Pixel = 97;
			11854: Pixel = 91;
			11855: Pixel = 89;
			11856: Pixel = 76;
			11857: Pixel = 74;
			11858: Pixel = 109;
			11859: Pixel = 142;
			11860: Pixel = 159;
			11861: Pixel = 173;
			11862: Pixel = 178;
			11863: Pixel = 179;
			11864: Pixel = 180;
			11865: Pixel = 177;
			11866: Pixel = 165;
			11867: Pixel = 143;
			11868: Pixel = 115;
			11869: Pixel = 84;
			11870: Pixel = 80;
			11871: Pixel = 90;
			11872: Pixel = 98;
			11873: Pixel = 102;
			11874: Pixel = 105;
			11875: Pixel = 104;
			11876: Pixel = 103;
			11877: Pixel = 108;
			11878: Pixel = 97;
			11879: Pixel = 65;
			11880: Pixel = 45;
			11881: Pixel = 104;
			11882: Pixel = 137;
			11883: Pixel = 176;
			11884: Pixel = 238;
			11885: Pixel = 169;
			11886: Pixel = 62;
			11887: Pixel = 36;
			11888: Pixel = 30;
			11889: Pixel = 54;
			11890: Pixel = 91;
			11891: Pixel = 67;
			11892: Pixel = 56;
			11893: Pixel = 73;
			11894: Pixel = 71;
			11895: Pixel = 74;
			11896: Pixel = 100;
			11897: Pixel = 102;
			11898: Pixel = 119;
			11899: Pixel = 53;
			11900: Pixel = 44;
			11901: Pixel = 52;
			11902: Pixel = 45;
			11903: Pixel = 51;
			11904: Pixel = 70;
			11905: Pixel = 49;
			11906: Pixel = 45;
			11907: Pixel = 47;
			11908: Pixel = 45;
			11909: Pixel = 38;
			11910: Pixel = 36;
			11911: Pixel = 86;
			11912: Pixel = 108;
			11913: Pixel = 149;
			11914: Pixel = 162;
			11915: Pixel = 175;
			11916: Pixel = 193;
			11917: Pixel = 202;
			11918: Pixel = 186;
			11919: Pixel = 120;
			11920: Pixel = 113;
			11921: Pixel = 129;
			11922: Pixel = 127;
			11923: Pixel = 92;
			11924: Pixel = 59;
			11925: Pixel = 110;
			11926: Pixel = 111;
			11927: Pixel = 81;
			11928: Pixel = 109;
			11929: Pixel = 192;
			11930: Pixel = 212;
			11931: Pixel = 197;
			11932: Pixel = 148;
			11933: Pixel = 111;
			11934: Pixel = 117;
			11935: Pixel = 115;
			11936: Pixel = 120;
			11937: Pixel = 128;
			11938: Pixel = 139;
			11939: Pixel = 161;
			11940: Pixel = 196;
			11941: Pixel = 225;
			11942: Pixel = 158;
			11943: Pixel = 103;
			11944: Pixel = 124;
			11945: Pixel = 91;
			11946: Pixel = 88;
			11947: Pixel = 124;
			11948: Pixel = 181;
			11949: Pixel = 129;
			11950: Pixel = 61;
			11951: Pixel = 45;
			11952: Pixel = 47;
			11953: Pixel = 47;
			11954: Pixel = 40;
			11955: Pixel = 60;
			11956: Pixel = 59;
			11957: Pixel = 124;
			11958: Pixel = 164;
			11959: Pixel = 79;
			11960: Pixel = 87;
			11961: Pixel = 65;
			11962: Pixel = 49;
			11963: Pixel = 50;
			11964: Pixel = 52;
			11965: Pixel = 55;
			11966: Pixel = 42;
			11967: Pixel = 60;
			11968: Pixel = 130;
			11969: Pixel = 141;
			11970: Pixel = 139;
			11971: Pixel = 156;
			11972: Pixel = 157;
			11973: Pixel = 155;
			11974: Pixel = 154;
			11975: Pixel = 153;
			11976: Pixel = 152;
			11977: Pixel = 151;
			11978: Pixel = 152;
			11979: Pixel = 152;
			11980: Pixel = 151;
			11981: Pixel = 152;
			11982: Pixel = 153;
			11983: Pixel = 152;
			11984: Pixel = 152;
			11985: Pixel = 151;
			11986: Pixel = 151;
			11987: Pixel = 148;
			11988: Pixel = 147;
			11989: Pixel = 146;
			11990: Pixel = 144;
			11991: Pixel = 143;
			11992: Pixel = 139;
			11993: Pixel = 136;
			11994: Pixel = 132;
			11995: Pixel = 128;
			11996: Pixel = 133;
			11997: Pixel = 143;
			11998: Pixel = 158;
			11999: Pixel = 172;
			12000: Pixel = 101;
			12001: Pixel = 100;
			12002: Pixel = 98;
			12003: Pixel = 97;
			12004: Pixel = 91;
			12005: Pixel = 88;
			12006: Pixel = 77;
			12007: Pixel = 74;
			12008: Pixel = 110;
			12009: Pixel = 142;
			12010: Pixel = 159;
			12011: Pixel = 172;
			12012: Pixel = 178;
			12013: Pixel = 179;
			12014: Pixel = 180;
			12015: Pixel = 179;
			12016: Pixel = 166;
			12017: Pixel = 146;
			12018: Pixel = 117;
			12019: Pixel = 87;
			12020: Pixel = 84;
			12021: Pixel = 93;
			12022: Pixel = 100;
			12023: Pixel = 107;
			12024: Pixel = 109;
			12025: Pixel = 111;
			12026: Pixel = 111;
			12027: Pixel = 55;
			12028: Pixel = 44;
			12029: Pixel = 93;
			12030: Pixel = 130;
			12031: Pixel = 157;
			12032: Pixel = 178;
			12033: Pixel = 198;
			12034: Pixel = 151;
			12035: Pixel = 60;
			12036: Pixel = 72;
			12037: Pixel = 54;
			12038: Pixel = 73;
			12039: Pixel = 107;
			12040: Pixel = 93;
			12041: Pixel = 44;
			12042: Pixel = 51;
			12043: Pixel = 76;
			12044: Pixel = 84;
			12045: Pixel = 78;
			12046: Pixel = 110;
			12047: Pixel = 97;
			12048: Pixel = 127;
			12049: Pixel = 81;
			12050: Pixel = 54;
			12051: Pixel = 48;
			12052: Pixel = 39;
			12053: Pixel = 45;
			12054: Pixel = 47;
			12055: Pixel = 54;
			12056: Pixel = 47;
			12057: Pixel = 50;
			12058: Pixel = 44;
			12059: Pixel = 30;
			12060: Pixel = 56;
			12061: Pixel = 123;
			12062: Pixel = 137;
			12063: Pixel = 182;
			12064: Pixel = 170;
			12065: Pixel = 192;
			12066: Pixel = 204;
			12067: Pixel = 183;
			12068: Pixel = 113;
			12069: Pixel = 118;
			12070: Pixel = 128;
			12071: Pixel = 132;
			12072: Pixel = 145;
			12073: Pixel = 135;
			12074: Pixel = 109;
			12075: Pixel = 102;
			12076: Pixel = 124;
			12077: Pixel = 134;
			12078: Pixel = 160;
			12079: Pixel = 180;
			12080: Pixel = 185;
			12081: Pixel = 177;
			12082: Pixel = 157;
			12083: Pixel = 139;
			12084: Pixel = 129;
			12085: Pixel = 122;
			12086: Pixel = 122;
			12087: Pixel = 129;
			12088: Pixel = 135;
			12089: Pixel = 161;
			12090: Pixel = 201;
			12091: Pixel = 224;
			12092: Pixel = 164;
			12093: Pixel = 112;
			12094: Pixel = 130;
			12095: Pixel = 136;
			12096: Pixel = 140;
			12097: Pixel = 172;
			12098: Pixel = 152;
			12099: Pixel = 97;
			12100: Pixel = 54;
			12101: Pixel = 63;
			12102: Pixel = 55;
			12103: Pixel = 52;
			12104: Pixel = 51;
			12105: Pixel = 65;
			12106: Pixel = 57;
			12107: Pixel = 114;
			12108: Pixel = 172;
			12109: Pixel = 87;
			12110: Pixel = 86;
			12111: Pixel = 64;
			12112: Pixel = 47;
			12113: Pixel = 46;
			12114: Pixel = 48;
			12115: Pixel = 54;
			12116: Pixel = 46;
			12117: Pixel = 84;
			12118: Pixel = 139;
			12119: Pixel = 135;
			12120: Pixel = 144;
			12121: Pixel = 159;
			12122: Pixel = 155;
			12123: Pixel = 155;
			12124: Pixel = 152;
			12125: Pixel = 152;
			12126: Pixel = 149;
			12127: Pixel = 150;
			12128: Pixel = 154;
			12129: Pixel = 162;
			12130: Pixel = 152;
			12131: Pixel = 152;
			12132: Pixel = 154;
			12133: Pixel = 153;
			12134: Pixel = 150;
			12135: Pixel = 149;
			12136: Pixel = 148;
			12137: Pixel = 146;
			12138: Pixel = 144;
			12139: Pixel = 144;
			12140: Pixel = 138;
			12141: Pixel = 138;
			12142: Pixel = 137;
			12143: Pixel = 131;
			12144: Pixel = 134;
			12145: Pixel = 149;
			12146: Pixel = 164;
			12147: Pixel = 175;
			12148: Pixel = 181;
			12149: Pixel = 187;
			12150: Pixel = 103;
			12151: Pixel = 103;
			12152: Pixel = 102;
			12153: Pixel = 97;
			12154: Pixel = 89;
			12155: Pixel = 85;
			12156: Pixel = 77;
			12157: Pixel = 72;
			12158: Pixel = 108;
			12159: Pixel = 143;
			12160: Pixel = 160;
			12161: Pixel = 172;
			12162: Pixel = 177;
			12163: Pixel = 180;
			12164: Pixel = 183;
			12165: Pixel = 181;
			12166: Pixel = 169;
			12167: Pixel = 148;
			12168: Pixel = 119;
			12169: Pixel = 86;
			12170: Pixel = 84;
			12171: Pixel = 96;
			12172: Pixel = 102;
			12173: Pixel = 109;
			12174: Pixel = 110;
			12175: Pixel = 115;
			12176: Pixel = 117;
			12177: Pixel = 45;
			12178: Pixel = 99;
			12179: Pixel = 152;
			12180: Pixel = 151;
			12181: Pixel = 132;
			12182: Pixel = 149;
			12183: Pixel = 108;
			12184: Pixel = 47;
			12185: Pixel = 41;
			12186: Pixel = 70;
			12187: Pixel = 121;
			12188: Pixel = 82;
			12189: Pixel = 88;
			12190: Pixel = 66;
			12191: Pixel = 31;
			12192: Pixel = 65;
			12193: Pixel = 79;
			12194: Pixel = 85;
			12195: Pixel = 61;
			12196: Pixel = 107;
			12197: Pixel = 121;
			12198: Pixel = 119;
			12199: Pixel = 103;
			12200: Pixel = 75;
			12201: Pixel = 39;
			12202: Pixel = 44;
			12203: Pixel = 44;
			12204: Pixel = 47;
			12205: Pixel = 45;
			12206: Pixel = 50;
			12207: Pixel = 48;
			12208: Pixel = 37;
			12209: Pixel = 28;
			12210: Pixel = 105;
			12211: Pixel = 116;
			12212: Pixel = 167;
			12213: Pixel = 172;
			12214: Pixel = 181;
			12215: Pixel = 203;
			12216: Pixel = 188;
			12217: Pixel = 105;
			12218: Pixel = 110;
			12219: Pixel = 133;
			12220: Pixel = 137;
			12221: Pixel = 138;
			12222: Pixel = 144;
			12223: Pixel = 144;
			12224: Pixel = 141;
			12225: Pixel = 136;
			12226: Pixel = 117;
			12227: Pixel = 110;
			12228: Pixel = 127;
			12229: Pixel = 125;
			12230: Pixel = 122;
			12231: Pixel = 153;
			12232: Pixel = 167;
			12233: Pixel = 155;
			12234: Pixel = 127;
			12235: Pixel = 123;
			12236: Pixel = 128;
			12237: Pixel = 127;
			12238: Pixel = 134;
			12239: Pixel = 156;
			12240: Pixel = 195;
			12241: Pixel = 225;
			12242: Pixel = 186;
			12243: Pixel = 157;
			12244: Pixel = 143;
			12245: Pixel = 133;
			12246: Pixel = 122;
			12247: Pixel = 118;
			12248: Pixel = 78;
			12249: Pixel = 68;
			12250: Pixel = 77;
			12251: Pixel = 79;
			12252: Pixel = 55;
			12253: Pixel = 48;
			12254: Pixel = 48;
			12255: Pixel = 70;
			12256: Pixel = 55;
			12257: Pixel = 106;
			12258: Pixel = 180;
			12259: Pixel = 99;
			12260: Pixel = 81;
			12261: Pixel = 59;
			12262: Pixel = 48;
			12263: Pixel = 47;
			12264: Pixel = 53;
			12265: Pixel = 53;
			12266: Pixel = 58;
			12267: Pixel = 114;
			12268: Pixel = 138;
			12269: Pixel = 133;
			12270: Pixel = 152;
			12271: Pixel = 159;
			12272: Pixel = 155;
			12273: Pixel = 154;
			12274: Pixel = 152;
			12275: Pixel = 152;
			12276: Pixel = 149;
			12277: Pixel = 149;
			12278: Pixel = 152;
			12279: Pixel = 155;
			12280: Pixel = 151;
			12281: Pixel = 151;
			12282: Pixel = 151;
			12283: Pixel = 153;
			12284: Pixel = 151;
			12285: Pixel = 147;
			12286: Pixel = 145;
			12287: Pixel = 143;
			12288: Pixel = 139;
			12289: Pixel = 138;
			12290: Pixel = 136;
			12291: Pixel = 134;
			12292: Pixel = 136;
			12293: Pixel = 147;
			12294: Pixel = 165;
			12295: Pixel = 178;
			12296: Pixel = 185;
			12297: Pixel = 188;
			12298: Pixel = 187;
			12299: Pixel = 188;
			12300: Pixel = 101;
			12301: Pixel = 101;
			12302: Pixel = 98;
			12303: Pixel = 94;
			12304: Pixel = 86;
			12305: Pixel = 84;
			12306: Pixel = 74;
			12307: Pixel = 69;
			12308: Pixel = 106;
			12309: Pixel = 141;
			12310: Pixel = 160;
			12311: Pixel = 173;
			12312: Pixel = 178;
			12313: Pixel = 180;
			12314: Pixel = 183;
			12315: Pixel = 182;
			12316: Pixel = 170;
			12317: Pixel = 149;
			12318: Pixel = 120;
			12319: Pixel = 85;
			12320: Pixel = 81;
			12321: Pixel = 93;
			12322: Pixel = 100;
			12323: Pixel = 107;
			12324: Pixel = 111;
			12325: Pixel = 105;
			12326: Pixel = 126;
			12327: Pixel = 138;
			12328: Pixel = 154;
			12329: Pixel = 149;
			12330: Pixel = 120;
			12331: Pixel = 73;
			12332: Pixel = 80;
			12333: Pixel = 76;
			12334: Pixel = 47;
			12335: Pixel = 48;
			12336: Pixel = 40;
			12337: Pixel = 90;
			12338: Pixel = 126;
			12339: Pixel = 127;
			12340: Pixel = 101;
			12341: Pixel = 57;
			12342: Pixel = 49;
			12343: Pixel = 74;
			12344: Pixel = 88;
			12345: Pixel = 87;
			12346: Pixel = 79;
			12347: Pixel = 107;
			12348: Pixel = 131;
			12349: Pixel = 117;
			12350: Pixel = 58;
			12351: Pixel = 49;
			12352: Pixel = 47;
			12353: Pixel = 48;
			12354: Pixel = 46;
			12355: Pixel = 48;
			12356: Pixel = 48;
			12357: Pixel = 45;
			12358: Pixel = 27;
			12359: Pixel = 67;
			12360: Pixel = 133;
			12361: Pixel = 131;
			12362: Pixel = 173;
			12363: Pixel = 172;
			12364: Pixel = 195;
			12365: Pixel = 197;
			12366: Pixel = 101;
			12367: Pixel = 94;
			12368: Pixel = 126;
			12369: Pixel = 135;
			12370: Pixel = 146;
			12371: Pixel = 148;
			12372: Pixel = 149;
			12373: Pixel = 147;
			12374: Pixel = 146;
			12375: Pixel = 145;
			12376: Pixel = 140;
			12377: Pixel = 135;
			12378: Pixel = 138;
			12379: Pixel = 141;
			12380: Pixel = 148;
			12381: Pixel = 158;
			12382: Pixel = 152;
			12383: Pixel = 153;
			12384: Pixel = 131;
			12385: Pixel = 128;
			12386: Pixel = 135;
			12387: Pixel = 127;
			12388: Pixel = 128;
			12389: Pixel = 152;
			12390: Pixel = 192;
			12391: Pixel = 223;
			12392: Pixel = 194;
			12393: Pixel = 161;
			12394: Pixel = 148;
			12395: Pixel = 134;
			12396: Pixel = 128;
			12397: Pixel = 123;
			12398: Pixel = 103;
			12399: Pixel = 94;
			12400: Pixel = 101;
			12401: Pixel = 83;
			12402: Pixel = 57;
			12403: Pixel = 44;
			12404: Pixel = 47;
			12405: Pixel = 67;
			12406: Pixel = 54;
			12407: Pixel = 102;
			12408: Pixel = 182;
			12409: Pixel = 110;
			12410: Pixel = 72;
			12411: Pixel = 56;
			12412: Pixel = 49;
			12413: Pixel = 45;
			12414: Pixel = 60;
			12415: Pixel = 45;
			12416: Pixel = 61;
			12417: Pixel = 130;
			12418: Pixel = 134;
			12419: Pixel = 135;
			12420: Pixel = 158;
			12421: Pixel = 157;
			12422: Pixel = 153;
			12423: Pixel = 154;
			12424: Pixel = 152;
			12425: Pixel = 150;
			12426: Pixel = 152;
			12427: Pixel = 151;
			12428: Pixel = 151;
			12429: Pixel = 149;
			12430: Pixel = 150;
			12431: Pixel = 150;
			12432: Pixel = 150;
			12433: Pixel = 150;
			12434: Pixel = 147;
			12435: Pixel = 146;
			12436: Pixel = 143;
			12437: Pixel = 141;
			12438: Pixel = 139;
			12439: Pixel = 135;
			12440: Pixel = 132;
			12441: Pixel = 137;
			12442: Pixel = 160;
			12443: Pixel = 178;
			12444: Pixel = 187;
			12445: Pixel = 190;
			12446: Pixel = 190;
			12447: Pixel = 189;
			12448: Pixel = 189;
			12449: Pixel = 188;
			12450: Pixel = 101;
			12451: Pixel = 95;
			12452: Pixel = 93;
			12453: Pixel = 87;
			12454: Pixel = 83;
			12455: Pixel = 81;
			12456: Pixel = 67;
			12457: Pixel = 60;
			12458: Pixel = 102;
			12459: Pixel = 140;
			12460: Pixel = 159;
			12461: Pixel = 171;
			12462: Pixel = 178;
			12463: Pixel = 181;
			12464: Pixel = 182;
			12465: Pixel = 182;
			12466: Pixel = 169;
			12467: Pixel = 150;
			12468: Pixel = 120;
			12469: Pixel = 84;
			12470: Pixel = 82;
			12471: Pixel = 93;
			12472: Pixel = 100;
			12473: Pixel = 108;
			12474: Pixel = 109;
			12475: Pixel = 107;
			12476: Pixel = 113;
			12477: Pixel = 149;
			12478: Pixel = 140;
			12479: Pixel = 113;
			12480: Pixel = 70;
			12481: Pixel = 69;
			12482: Pixel = 89;
			12483: Pixel = 58;
			12484: Pixel = 41;
			12485: Pixel = 66;
			12486: Pixel = 65;
			12487: Pixel = 86;
			12488: Pixel = 101;
			12489: Pixel = 92;
			12490: Pixel = 91;
			12491: Pixel = 43;
			12492: Pixel = 44;
			12493: Pixel = 72;
			12494: Pixel = 61;
			12495: Pixel = 102;
			12496: Pixel = 116;
			12497: Pixel = 90;
			12498: Pixel = 90;
			12499: Pixel = 100;
			12500: Pixel = 68;
			12501: Pixel = 47;
			12502: Pixel = 45;
			12503: Pixel = 45;
			12504: Pixel = 44;
			12505: Pixel = 51;
			12506: Pixel = 48;
			12507: Pixel = 43;
			12508: Pixel = 37;
			12509: Pixel = 120;
			12510: Pixel = 115;
			12511: Pixel = 163;
			12512: Pixel = 181;
			12513: Pixel = 190;
			12514: Pixel = 207;
			12515: Pixel = 107;
			12516: Pixel = 84;
			12517: Pixel = 116;
			12518: Pixel = 125;
			12519: Pixel = 136;
			12520: Pixel = 148;
			12521: Pixel = 154;
			12522: Pixel = 156;
			12523: Pixel = 162;
			12524: Pixel = 160;
			12525: Pixel = 157;
			12526: Pixel = 154;
			12527: Pixel = 155;
			12528: Pixel = 159;
			12529: Pixel = 166;
			12530: Pixel = 168;
			12531: Pixel = 166;
			12532: Pixel = 167;
			12533: Pixel = 157;
			12534: Pixel = 133;
			12535: Pixel = 138;
			12536: Pixel = 135;
			12537: Pixel = 128;
			12538: Pixel = 128;
			12539: Pixel = 150;
			12540: Pixel = 189;
			12541: Pixel = 221;
			12542: Pixel = 201;
			12543: Pixel = 179;
			12544: Pixel = 161;
			12545: Pixel = 153;
			12546: Pixel = 142;
			12547: Pixel = 130;
			12548: Pixel = 124;
			12549: Pixel = 114;
			12550: Pixel = 113;
			12551: Pixel = 92;
			12552: Pixel = 62;
			12553: Pixel = 48;
			12554: Pixel = 51;
			12555: Pixel = 67;
			12556: Pixel = 51;
			12557: Pixel = 98;
			12558: Pixel = 182;
			12559: Pixel = 116;
			12560: Pixel = 69;
			12561: Pixel = 55;
			12562: Pixel = 49;
			12563: Pixel = 45;
			12564: Pixel = 54;
			12565: Pixel = 39;
			12566: Pixel = 76;
			12567: Pixel = 137;
			12568: Pixel = 133;
			12569: Pixel = 142;
			12570: Pixel = 157;
			12571: Pixel = 155;
			12572: Pixel = 154;
			12573: Pixel = 152;
			12574: Pixel = 151;
			12575: Pixel = 149;
			12576: Pixel = 150;
			12577: Pixel = 151;
			12578: Pixel = 151;
			12579: Pixel = 149;
			12580: Pixel = 149;
			12581: Pixel = 149;
			12582: Pixel = 148;
			12583: Pixel = 148;
			12584: Pixel = 145;
			12585: Pixel = 144;
			12586: Pixel = 141;
			12587: Pixel = 141;
			12588: Pixel = 136;
			12589: Pixel = 129;
			12590: Pixel = 140;
			12591: Pixel = 170;
			12592: Pixel = 189;
			12593: Pixel = 193;
			12594: Pixel = 193;
			12595: Pixel = 192;
			12596: Pixel = 190;
			12597: Pixel = 189;
			12598: Pixel = 189;
			12599: Pixel = 189;
			12600: Pixel = 94;
			12601: Pixel = 91;
			12602: Pixel = 88;
			12603: Pixel = 84;
			12604: Pixel = 80;
			12605: Pixel = 77;
			12606: Pixel = 64;
			12607: Pixel = 62;
			12608: Pixel = 98;
			12609: Pixel = 139;
			12610: Pixel = 158;
			12611: Pixel = 171;
			12612: Pixel = 178;
			12613: Pixel = 180;
			12614: Pixel = 182;
			12615: Pixel = 181;
			12616: Pixel = 169;
			12617: Pixel = 149;
			12618: Pixel = 120;
			12619: Pixel = 86;
			12620: Pixel = 81;
			12621: Pixel = 92;
			12622: Pixel = 99;
			12623: Pixel = 105;
			12624: Pixel = 107;
			12625: Pixel = 109;
			12626: Pixel = 118;
			12627: Pixel = 114;
			12628: Pixel = 130;
			12629: Pixel = 125;
			12630: Pixel = 123;
			12631: Pixel = 120;
			12632: Pixel = 67;
			12633: Pixel = 51;
			12634: Pixel = 58;
			12635: Pixel = 86;
			12636: Pixel = 101;
			12637: Pixel = 118;
			12638: Pixel = 74;
			12639: Pixel = 95;
			12640: Pixel = 64;
			12641: Pixel = 34;
			12642: Pixel = 47;
			12643: Pixel = 88;
			12644: Pixel = 95;
			12645: Pixel = 71;
			12646: Pixel = 114;
			12647: Pixel = 101;
			12648: Pixel = 118;
			12649: Pixel = 122;
			12650: Pixel = 52;
			12651: Pixel = 52;
			12652: Pixel = 49;
			12653: Pixel = 48;
			12654: Pixel = 43;
			12655: Pixel = 47;
			12656: Pixel = 51;
			12657: Pixel = 39;
			12658: Pixel = 84;
			12659: Pixel = 128;
			12660: Pixel = 128;
			12661: Pixel = 181;
			12662: Pixel = 185;
			12663: Pixel = 209;
			12664: Pixel = 124;
			12665: Pixel = 63;
			12666: Pixel = 108;
			12667: Pixel = 119;
			12668: Pixel = 126;
			12669: Pixel = 136;
			12670: Pixel = 145;
			12671: Pixel = 153;
			12672: Pixel = 160;
			12673: Pixel = 167;
			12674: Pixel = 165;
			12675: Pixel = 174;
			12676: Pixel = 170;
			12677: Pixel = 168;
			12678: Pixel = 171;
			12679: Pixel = 172;
			12680: Pixel = 169;
			12681: Pixel = 170;
			12682: Pixel = 165;
			12683: Pixel = 150;
			12684: Pixel = 138;
			12685: Pixel = 142;
			12686: Pixel = 132;
			12687: Pixel = 129;
			12688: Pixel = 126;
			12689: Pixel = 144;
			12690: Pixel = 185;
			12691: Pixel = 219;
			12692: Pixel = 206;
			12693: Pixel = 180;
			12694: Pixel = 169;
			12695: Pixel = 154;
			12696: Pixel = 145;
			12697: Pixel = 136;
			12698: Pixel = 130;
			12699: Pixel = 122;
			12700: Pixel = 117;
			12701: Pixel = 97;
			12702: Pixel = 62;
			12703: Pixel = 48;
			12704: Pixel = 53;
			12705: Pixel = 68;
			12706: Pixel = 46;
			12707: Pixel = 89;
			12708: Pixel = 185;
			12709: Pixel = 127;
			12710: Pixel = 60;
			12711: Pixel = 50;
			12712: Pixel = 50;
			12713: Pixel = 46;
			12714: Pixel = 50;
			12715: Pixel = 42;
			12716: Pixel = 98;
			12717: Pixel = 139;
			12718: Pixel = 132;
			12719: Pixel = 150;
			12720: Pixel = 159;
			12721: Pixel = 155;
			12722: Pixel = 154;
			12723: Pixel = 151;
			12724: Pixel = 151;
			12725: Pixel = 151;
			12726: Pixel = 150;
			12727: Pixel = 152;
			12728: Pixel = 151;
			12729: Pixel = 148;
			12730: Pixel = 149;
			12731: Pixel = 148;
			12732: Pixel = 146;
			12733: Pixel = 145;
			12734: Pixel = 144;
			12735: Pixel = 141;
			12736: Pixel = 139;
			12737: Pixel = 137;
			12738: Pixel = 130;
			12739: Pixel = 140;
			12740: Pixel = 173;
			12741: Pixel = 191;
			12742: Pixel = 197;
			12743: Pixel = 197;
			12744: Pixel = 193;
			12745: Pixel = 191;
			12746: Pixel = 189;
			12747: Pixel = 188;
			12748: Pixel = 189;
			12749: Pixel = 190;
			12750: Pixel = 90;
			12751: Pixel = 94;
			12752: Pixel = 85;
			12753: Pixel = 83;
			12754: Pixel = 79;
			12755: Pixel = 74;
			12756: Pixel = 63;
			12757: Pixel = 60;
			12758: Pixel = 100;
			12759: Pixel = 137;
			12760: Pixel = 159;
			12761: Pixel = 171;
			12762: Pixel = 176;
			12763: Pixel = 179;
			12764: Pixel = 181;
			12765: Pixel = 180;
			12766: Pixel = 169;
			12767: Pixel = 150;
			12768: Pixel = 119;
			12769: Pixel = 83;
			12770: Pixel = 80;
			12771: Pixel = 90;
			12772: Pixel = 96;
			12773: Pixel = 105;
			12774: Pixel = 126;
			12775: Pixel = 140;
			12776: Pixel = 144;
			12777: Pixel = 147;
			12778: Pixel = 149;
			12779: Pixel = 103;
			12780: Pixel = 97;
			12781: Pixel = 76;
			12782: Pixel = 59;
			12783: Pixel = 62;
			12784: Pixel = 74;
			12785: Pixel = 92;
			12786: Pixel = 97;
			12787: Pixel = 104;
			12788: Pixel = 120;
			12789: Pixel = 86;
			12790: Pixel = 41;
			12791: Pixel = 41;
			12792: Pixel = 44;
			12793: Pixel = 52;
			12794: Pixel = 88;
			12795: Pixel = 102;
			12796: Pixel = 108;
			12797: Pixel = 111;
			12798: Pixel = 97;
			12799: Pixel = 81;
			12800: Pixel = 119;
			12801: Pixel = 87;
			12802: Pixel = 48;
			12803: Pixel = 48;
			12804: Pixel = 46;
			12805: Pixel = 46;
			12806: Pixel = 44;
			12807: Pixel = 42;
			12808: Pixel = 129;
			12809: Pixel = 112;
			12810: Pixel = 163;
			12811: Pixel = 186;
			12812: Pixel = 208;
			12813: Pixel = 151;
			12814: Pixel = 44;
			12815: Pixel = 84;
			12816: Pixel = 111;
			12817: Pixel = 121;
			12818: Pixel = 127;
			12819: Pixel = 135;
			12820: Pixel = 144;
			12821: Pixel = 152;
			12822: Pixel = 157;
			12823: Pixel = 167;
			12824: Pixel = 170;
			12825: Pixel = 175;
			12826: Pixel = 174;
			12827: Pixel = 175;
			12828: Pixel = 175;
			12829: Pixel = 171;
			12830: Pixel = 175;
			12831: Pixel = 175;
			12832: Pixel = 163;
			12833: Pixel = 151;
			12834: Pixel = 144;
			12835: Pixel = 144;
			12836: Pixel = 134;
			12837: Pixel = 130;
			12838: Pixel = 127;
			12839: Pixel = 138;
			12840: Pixel = 178;
			12841: Pixel = 218;
			12842: Pixel = 211;
			12843: Pixel = 178;
			12844: Pixel = 169;
			12845: Pixel = 158;
			12846: Pixel = 144;
			12847: Pixel = 135;
			12848: Pixel = 132;
			12849: Pixel = 127;
			12850: Pixel = 122;
			12851: Pixel = 103;
			12852: Pixel = 61;
			12853: Pixel = 50;
			12854: Pixel = 58;
			12855: Pixel = 69;
			12856: Pixel = 45;
			12857: Pixel = 82;
			12858: Pixel = 179;
			12859: Pixel = 138;
			12860: Pixel = 57;
			12861: Pixel = 46;
			12862: Pixel = 49;
			12863: Pixel = 50;
			12864: Pixel = 47;
			12865: Pixel = 52;
			12866: Pixel = 121;
			12867: Pixel = 139;
			12868: Pixel = 135;
			12869: Pixel = 157;
			12870: Pixel = 158;
			12871: Pixel = 154;
			12872: Pixel = 153;
			12873: Pixel = 153;
			12874: Pixel = 151;
			12875: Pixel = 151;
			12876: Pixel = 151;
			12877: Pixel = 151;
			12878: Pixel = 151;
			12879: Pixel = 148;
			12880: Pixel = 147;
			12881: Pixel = 145;
			12882: Pixel = 146;
			12883: Pixel = 145;
			12884: Pixel = 142;
			12885: Pixel = 138;
			12886: Pixel = 137;
			12887: Pixel = 132;
			12888: Pixel = 138;
			12889: Pixel = 170;
			12890: Pixel = 190;
			12891: Pixel = 197;
			12892: Pixel = 197;
			12893: Pixel = 196;
			12894: Pixel = 193;
			12895: Pixel = 191;
			12896: Pixel = 189;
			12897: Pixel = 190;
			12898: Pixel = 192;
			12899: Pixel = 193;
			12900: Pixel = 84;
			12901: Pixel = 86;
			12902: Pixel = 80;
			12903: Pixel = 79;
			12904: Pixel = 79;
			12905: Pixel = 72;
			12906: Pixel = 63;
			12907: Pixel = 58;
			12908: Pixel = 100;
			12909: Pixel = 138;
			12910: Pixel = 158;
			12911: Pixel = 172;
			12912: Pixel = 176;
			12913: Pixel = 178;
			12914: Pixel = 181;
			12915: Pixel = 180;
			12916: Pixel = 168;
			12917: Pixel = 149;
			12918: Pixel = 119;
			12919: Pixel = 83;
			12920: Pixel = 79;
			12921: Pixel = 88;
			12922: Pixel = 103;
			12923: Pixel = 122;
			12924: Pixel = 124;
			12925: Pixel = 128;
			12926: Pixel = 128;
			12927: Pixel = 116;
			12928: Pixel = 82;
			12929: Pixel = 63;
			12930: Pixel = 75;
			12931: Pixel = 60;
			12932: Pixel = 56;
			12933: Pixel = 71;
			12934: Pixel = 86;
			12935: Pixel = 84;
			12936: Pixel = 119;
			12937: Pixel = 120;
			12938: Pixel = 95;
			12939: Pixel = 48;
			12940: Pixel = 50;
			12941: Pixel = 46;
			12942: Pixel = 44;
			12943: Pixel = 46;
			12944: Pixel = 54;
			12945: Pixel = 74;
			12946: Pixel = 84;
			12947: Pixel = 65;
			12948: Pixel = 21;
			12949: Pixel = 87;
			12950: Pixel = 142;
			12951: Pixel = 92;
			12952: Pixel = 51;
			12953: Pixel = 45;
			12954: Pixel = 46;
			12955: Pixel = 47;
			12956: Pixel = 35;
			12957: Pixel = 86;
			12958: Pixel = 132;
			12959: Pixel = 131;
			12960: Pixel = 183;
			12961: Pixel = 196;
			12962: Pixel = 187;
			12963: Pixel = 50;
			12964: Pixel = 51;
			12965: Pixel = 95;
			12966: Pixel = 116;
			12967: Pixel = 123;
			12968: Pixel = 125;
			12969: Pixel = 134;
			12970: Pixel = 143;
			12971: Pixel = 150;
			12972: Pixel = 156;
			12973: Pixel = 165;
			12974: Pixel = 172;
			12975: Pixel = 176;
			12976: Pixel = 178;
			12977: Pixel = 177;
			12978: Pixel = 176;
			12979: Pixel = 176;
			12980: Pixel = 176;
			12981: Pixel = 170;
			12982: Pixel = 162;
			12983: Pixel = 153;
			12984: Pixel = 148;
			12985: Pixel = 145;
			12986: Pixel = 137;
			12987: Pixel = 132;
			12988: Pixel = 128;
			12989: Pixel = 136;
			12990: Pixel = 174;
			12991: Pixel = 217;
			12992: Pixel = 215;
			12993: Pixel = 179;
			12994: Pixel = 162;
			12995: Pixel = 160;
			12996: Pixel = 149;
			12997: Pixel = 137;
			12998: Pixel = 132;
			12999: Pixel = 128;
			13000: Pixel = 125;
			13001: Pixel = 100;
			13002: Pixel = 57;
			13003: Pixel = 52;
			13004: Pixel = 57;
			13005: Pixel = 73;
			13006: Pixel = 46;
			13007: Pixel = 75;
			13008: Pixel = 167;
			13009: Pixel = 149;
			13010: Pixel = 65;
			13011: Pixel = 38;
			13012: Pixel = 48;
			13013: Pixel = 52;
			13014: Pixel = 41;
			13015: Pixel = 64;
			13016: Pixel = 134;
			13017: Pixel = 137;
			13018: Pixel = 142;
			13019: Pixel = 160;
			13020: Pixel = 157;
			13021: Pixel = 154;
			13022: Pixel = 154;
			13023: Pixel = 153;
			13024: Pixel = 150;
			13025: Pixel = 152;
			13026: Pixel = 150;
			13027: Pixel = 149;
			13028: Pixel = 149;
			13029: Pixel = 148;
			13030: Pixel = 146;
			13031: Pixel = 145;
			13032: Pixel = 145;
			13033: Pixel = 143;
			13034: Pixel = 142;
			13035: Pixel = 137;
			13036: Pixel = 132;
			13037: Pixel = 132;
			13038: Pixel = 162;
			13039: Pixel = 188;
			13040: Pixel = 194;
			13041: Pixel = 194;
			13042: Pixel = 194;
			13043: Pixel = 195;
			13044: Pixel = 194;
			13045: Pixel = 192;
			13046: Pixel = 191;
			13047: Pixel = 194;
			13048: Pixel = 198;
			13049: Pixel = 200;
			13050: Pixel = 82;
			13051: Pixel = 78;
			13052: Pixel = 77;
			13053: Pixel = 75;
			13054: Pixel = 74;
			13055: Pixel = 71;
			13056: Pixel = 62;
			13057: Pixel = 58;
			13058: Pixel = 97;
			13059: Pixel = 138;
			13060: Pixel = 157;
			13061: Pixel = 170;
			13062: Pixel = 176;
			13063: Pixel = 179;
			13064: Pixel = 179;
			13065: Pixel = 178;
			13066: Pixel = 167;
			13067: Pixel = 149;
			13068: Pixel = 120;
			13069: Pixel = 84;
			13070: Pixel = 81;
			13071: Pixel = 91;
			13072: Pixel = 101;
			13073: Pixel = 106;
			13074: Pixel = 107;
			13075: Pixel = 121;
			13076: Pixel = 104;
			13077: Pixel = 76;
			13078: Pixel = 96;
			13079: Pixel = 98;
			13080: Pixel = 89;
			13081: Pixel = 68;
			13082: Pixel = 70;
			13083: Pixel = 106;
			13084: Pixel = 61;
			13085: Pixel = 94;
			13086: Pixel = 131;
			13087: Pixel = 80;
			13088: Pixel = 70;
			13089: Pixel = 56;
			13090: Pixel = 43;
			13091: Pixel = 50;
			13092: Pixel = 49;
			13093: Pixel = 50;
			13094: Pixel = 49;
			13095: Pixel = 56;
			13096: Pixel = 58;
			13097: Pixel = 62;
			13098: Pixel = 33;
			13099: Pixel = 89;
			13100: Pixel = 133;
			13101: Pixel = 127;
			13102: Pixel = 50;
			13103: Pixel = 37;
			13104: Pixel = 40;
			13105: Pixel = 38;
			13106: Pixel = 38;
			13107: Pixel = 127;
			13108: Pixel = 117;
			13109: Pixel = 171;
			13110: Pixel = 192;
			13111: Pixel = 201;
			13112: Pixel = 88;
			13113: Pixel = 34;
			13114: Pixel = 64;
			13115: Pixel = 98;
			13116: Pixel = 118;
			13117: Pixel = 123;
			13118: Pixel = 127;
			13119: Pixel = 131;
			13120: Pixel = 138;
			13121: Pixel = 147;
			13122: Pixel = 149;
			13123: Pixel = 160;
			13124: Pixel = 169;
			13125: Pixel = 174;
			13126: Pixel = 178;
			13127: Pixel = 181;
			13128: Pixel = 177;
			13129: Pixel = 172;
			13130: Pixel = 172;
			13131: Pixel = 167;
			13132: Pixel = 158;
			13133: Pixel = 149;
			13134: Pixel = 146;
			13135: Pixel = 145;
			13136: Pixel = 137;
			13137: Pixel = 128;
			13138: Pixel = 129;
			13139: Pixel = 137;
			13140: Pixel = 168;
			13141: Pixel = 215;
			13142: Pixel = 219;
			13143: Pixel = 180;
			13144: Pixel = 164;
			13145: Pixel = 160;
			13146: Pixel = 150;
			13147: Pixel = 141;
			13148: Pixel = 133;
			13149: Pixel = 129;
			13150: Pixel = 125;
			13151: Pixel = 92;
			13152: Pixel = 55;
			13153: Pixel = 51;
			13154: Pixel = 52;
			13155: Pixel = 76;
			13156: Pixel = 42;
			13157: Pixel = 69;
			13158: Pixel = 162;
			13159: Pixel = 153;
			13160: Pixel = 76;
			13161: Pixel = 33;
			13162: Pixel = 57;
			13163: Pixel = 54;
			13164: Pixel = 41;
			13165: Pixel = 84;
			13166: Pixel = 140;
			13167: Pixel = 137;
			13168: Pixel = 152;
			13169: Pixel = 162;
			13170: Pixel = 156;
			13171: Pixel = 152;
			13172: Pixel = 154;
			13173: Pixel = 153;
			13174: Pixel = 150;
			13175: Pixel = 149;
			13176: Pixel = 149;
			13177: Pixel = 148;
			13178: Pixel = 147;
			13179: Pixel = 147;
			13180: Pixel = 147;
			13181: Pixel = 144;
			13182: Pixel = 145;
			13183: Pixel = 142;
			13184: Pixel = 139;
			13185: Pixel = 135;
			13186: Pixel = 126;
			13187: Pixel = 148;
			13188: Pixel = 183;
			13189: Pixel = 194;
			13190: Pixel = 195;
			13191: Pixel = 192;
			13192: Pixel = 193;
			13193: Pixel = 194;
			13194: Pixel = 194;
			13195: Pixel = 194;
			13196: Pixel = 196;
			13197: Pixel = 201;
			13198: Pixel = 203;
			13199: Pixel = 203;
			13200: Pixel = 77;
			13201: Pixel = 75;
			13202: Pixel = 74;
			13203: Pixel = 75;
			13204: Pixel = 70;
			13205: Pixel = 68;
			13206: Pixel = 59;
			13207: Pixel = 57;
			13208: Pixel = 94;
			13209: Pixel = 139;
			13210: Pixel = 156;
			13211: Pixel = 169;
			13212: Pixel = 174;
			13213: Pixel = 174;
			13214: Pixel = 175;
			13215: Pixel = 175;
			13216: Pixel = 167;
			13217: Pixel = 150;
			13218: Pixel = 121;
			13219: Pixel = 82;
			13220: Pixel = 80;
			13221: Pixel = 93;
			13222: Pixel = 99;
			13223: Pixel = 104;
			13224: Pixel = 105;
			13225: Pixel = 113;
			13226: Pixel = 102;
			13227: Pixel = 128;
			13228: Pixel = 113;
			13229: Pixel = 82;
			13230: Pixel = 100;
			13231: Pixel = 87;
			13232: Pixel = 106;
			13233: Pixel = 65;
			13234: Pixel = 53;
			13235: Pixel = 68;
			13236: Pixel = 117;
			13237: Pixel = 95;
			13238: Pixel = 62;
			13239: Pixel = 55;
			13240: Pixel = 49;
			13241: Pixel = 54;
			13242: Pixel = 49;
			13243: Pixel = 48;
			13244: Pixel = 46;
			13245: Pixel = 61;
			13246: Pixel = 55;
			13247: Pixel = 53;
			13248: Pixel = 39;
			13249: Pixel = 92;
			13250: Pixel = 103;
			13251: Pixel = 146;
			13252: Pixel = 110;
			13253: Pixel = 35;
			13254: Pixel = 38;
			13255: Pixel = 30;
			13256: Pixel = 78;
			13257: Pixel = 127;
			13258: Pixel = 127;
			13259: Pixel = 189;
			13260: Pixel = 211;
			13261: Pixel = 142;
			13262: Pixel = 32;
			13263: Pixel = 54;
			13264: Pixel = 61;
			13265: Pixel = 96;
			13266: Pixel = 117;
			13267: Pixel = 123;
			13268: Pixel = 129;
			13269: Pixel = 133;
			13270: Pixel = 139;
			13271: Pixel = 145;
			13272: Pixel = 150;
			13273: Pixel = 154;
			13274: Pixel = 160;
			13275: Pixel = 169;
			13276: Pixel = 175;
			13277: Pixel = 176;
			13278: Pixel = 177;
			13279: Pixel = 171;
			13280: Pixel = 170;
			13281: Pixel = 163;
			13282: Pixel = 156;
			13283: Pixel = 145;
			13284: Pixel = 139;
			13285: Pixel = 140;
			13286: Pixel = 134;
			13287: Pixel = 125;
			13288: Pixel = 127;
			13289: Pixel = 139;
			13290: Pixel = 161;
			13291: Pixel = 204;
			13292: Pixel = 222;
			13293: Pixel = 181;
			13294: Pixel = 161;
			13295: Pixel = 157;
			13296: Pixel = 149;
			13297: Pixel = 143;
			13298: Pixel = 134;
			13299: Pixel = 129;
			13300: Pixel = 122;
			13301: Pixel = 84;
			13302: Pixel = 49;
			13303: Pixel = 48;
			13304: Pixel = 52;
			13305: Pixel = 76;
			13306: Pixel = 40;
			13307: Pixel = 60;
			13308: Pixel = 164;
			13309: Pixel = 157;
			13310: Pixel = 95;
			13311: Pixel = 33;
			13312: Pixel = 55;
			13313: Pixel = 56;
			13314: Pixel = 47;
			13315: Pixel = 108;
			13316: Pixel = 141;
			13317: Pixel = 137;
			13318: Pixel = 166;
			13319: Pixel = 162;
			13320: Pixel = 154;
			13321: Pixel = 154;
			13322: Pixel = 154;
			13323: Pixel = 152;
			13324: Pixel = 151;
			13325: Pixel = 149;
			13326: Pixel = 147;
			13327: Pixel = 146;
			13328: Pixel = 147;
			13329: Pixel = 145;
			13330: Pixel = 143;
			13331: Pixel = 143;
			13332: Pixel = 143;
			13333: Pixel = 141;
			13334: Pixel = 136;
			13335: Pixel = 130;
			13336: Pixel = 135;
			13337: Pixel = 172;
			13338: Pixel = 193;
			13339: Pixel = 195;
			13340: Pixel = 194;
			13341: Pixel = 192;
			13342: Pixel = 193;
			13343: Pixel = 194;
			13344: Pixel = 196;
			13345: Pixel = 200;
			13346: Pixel = 204;
			13347: Pixel = 204;
			13348: Pixel = 205;
			13349: Pixel = 203;
			13350: Pixel = 77;
			13351: Pixel = 75;
			13352: Pixel = 74;
			13353: Pixel = 76;
			13354: Pixel = 71;
			13355: Pixel = 66;
			13356: Pixel = 55;
			13357: Pixel = 53;
			13358: Pixel = 96;
			13359: Pixel = 138;
			13360: Pixel = 156;
			13361: Pixel = 169;
			13362: Pixel = 174;
			13363: Pixel = 171;
			13364: Pixel = 176;
			13365: Pixel = 176;
			13366: Pixel = 164;
			13367: Pixel = 148;
			13368: Pixel = 121;
			13369: Pixel = 80;
			13370: Pixel = 72;
			13371: Pixel = 115;
			13372: Pixel = 103;
			13373: Pixel = 97;
			13374: Pixel = 127;
			13375: Pixel = 145;
			13376: Pixel = 128;
			13377: Pixel = 73;
			13378: Pixel = 67;
			13379: Pixel = 129;
			13380: Pixel = 98;
			13381: Pixel = 98;
			13382: Pixel = 52;
			13383: Pixel = 75;
			13384: Pixel = 77;
			13385: Pixel = 72;
			13386: Pixel = 130;
			13387: Pixel = 114;
			13388: Pixel = 71;
			13389: Pixel = 54;
			13390: Pixel = 62;
			13391: Pixel = 54;
			13392: Pixel = 42;
			13393: Pixel = 43;
			13394: Pixel = 40;
			13395: Pixel = 63;
			13396: Pixel = 70;
			13397: Pixel = 56;
			13398: Pixel = 53;
			13399: Pixel = 105;
			13400: Pixel = 131;
			13401: Pixel = 80;
			13402: Pixel = 155;
			13403: Pixel = 85;
			13404: Pixel = 29;
			13405: Pixel = 37;
			13406: Pixel = 117;
			13407: Pixel = 114;
			13408: Pixel = 163;
			13409: Pixel = 210;
			13410: Pixel = 194;
			13411: Pixel = 50;
			13412: Pixel = 37;
			13413: Pixel = 62;
			13414: Pixel = 60;
			13415: Pixel = 92;
			13416: Pixel = 111;
			13417: Pixel = 123;
			13418: Pixel = 128;
			13419: Pixel = 132;
			13420: Pixel = 137;
			13421: Pixel = 144;
			13422: Pixel = 151;
			13423: Pixel = 155;
			13424: Pixel = 159;
			13425: Pixel = 164;
			13426: Pixel = 172;
			13427: Pixel = 172;
			13428: Pixel = 172;
			13429: Pixel = 170;
			13430: Pixel = 167;
			13431: Pixel = 162;
			13432: Pixel = 154;
			13433: Pixel = 142;
			13434: Pixel = 133;
			13435: Pixel = 135;
			13436: Pixel = 131;
			13437: Pixel = 124;
			13438: Pixel = 124;
			13439: Pixel = 134;
			13440: Pixel = 155;
			13441: Pixel = 198;
			13442: Pixel = 224;
			13443: Pixel = 185;
			13444: Pixel = 158;
			13445: Pixel = 156;
			13446: Pixel = 148;
			13447: Pixel = 141;
			13448: Pixel = 134;
			13449: Pixel = 129;
			13450: Pixel = 118;
			13451: Pixel = 73;
			13452: Pixel = 44;
			13453: Pixel = 54;
			13454: Pixel = 58;
			13455: Pixel = 78;
			13456: Pixel = 41;
			13457: Pixel = 52;
			13458: Pixel = 154;
			13459: Pixel = 152;
			13460: Pixel = 111;
			13461: Pixel = 40;
			13462: Pixel = 53;
			13463: Pixel = 48;
			13464: Pixel = 56;
			13465: Pixel = 127;
			13466: Pixel = 139;
			13467: Pixel = 143;
			13468: Pixel = 162;
			13469: Pixel = 159;
			13470: Pixel = 156;
			13471: Pixel = 155;
			13472: Pixel = 153;
			13473: Pixel = 152;
			13474: Pixel = 151;
			13475: Pixel = 149;
			13476: Pixel = 148;
			13477: Pixel = 145;
			13478: Pixel = 145;
			13479: Pixel = 144;
			13480: Pixel = 144;
			13481: Pixel = 143;
			13482: Pixel = 141;
			13483: Pixel = 139;
			13484: Pixel = 134;
			13485: Pixel = 129;
			13486: Pixel = 156;
			13487: Pixel = 188;
			13488: Pixel = 195;
			13489: Pixel = 194;
			13490: Pixel = 192;
			13491: Pixel = 192;
			13492: Pixel = 193;
			13493: Pixel = 196;
			13494: Pixel = 201;
			13495: Pixel = 206;
			13496: Pixel = 208;
			13497: Pixel = 206;
			13498: Pixel = 202;
			13499: Pixel = 201;
			13500: Pixel = 78;
			13501: Pixel = 76;
			13502: Pixel = 77;
			13503: Pixel = 75;
			13504: Pixel = 69;
			13505: Pixel = 64;
			13506: Pixel = 54;
			13507: Pixel = 51;
			13508: Pixel = 96;
			13509: Pixel = 137;
			13510: Pixel = 155;
			13511: Pixel = 169;
			13512: Pixel = 172;
			13513: Pixel = 171;
			13514: Pixel = 175;
			13515: Pixel = 176;
			13516: Pixel = 164;
			13517: Pixel = 148;
			13518: Pixel = 118;
			13519: Pixel = 79;
			13520: Pixel = 69;
			13521: Pixel = 110;
			13522: Pixel = 125;
			13523: Pixel = 129;
			13524: Pixel = 136;
			13525: Pixel = 132;
			13526: Pixel = 86;
			13527: Pixel = 50;
			13528: Pixel = 120;
			13529: Pixel = 112;
			13530: Pixel = 96;
			13531: Pixel = 67;
			13532: Pixel = 57;
			13533: Pixel = 98;
			13534: Pixel = 92;
			13535: Pixel = 102;
			13536: Pixel = 128;
			13537: Pixel = 111;
			13538: Pixel = 99;
			13539: Pixel = 53;
			13540: Pixel = 61;
			13541: Pixel = 52;
			13542: Pixel = 37;
			13543: Pixel = 37;
			13544: Pixel = 46;
			13545: Pixel = 88;
			13546: Pixel = 99;
			13547: Pixel = 54;
			13548: Pixel = 82;
			13549: Pixel = 139;
			13550: Pixel = 192;
			13551: Pixel = 79;
			13552: Pixel = 90;
			13553: Pixel = 83;
			13554: Pixel = 16;
			13555: Pixel = 65;
			13556: Pixel = 133;
			13557: Pixel = 117;
			13558: Pixel = 194;
			13559: Pixel = 213;
			13560: Pixel = 88;
			13561: Pixel = 25;
			13562: Pixel = 43;
			13563: Pixel = 69;
			13564: Pixel = 60;
			13565: Pixel = 90;
			13566: Pixel = 110;
			13567: Pixel = 122;
			13568: Pixel = 128;
			13569: Pixel = 130;
			13570: Pixel = 135;
			13571: Pixel = 141;
			13572: Pixel = 149;
			13573: Pixel = 153;
			13574: Pixel = 158;
			13575: Pixel = 160;
			13576: Pixel = 163;
			13577: Pixel = 167;
			13578: Pixel = 168;
			13579: Pixel = 168;
			13580: Pixel = 165;
			13581: Pixel = 162;
			13582: Pixel = 152;
			13583: Pixel = 139;
			13584: Pixel = 132;
			13585: Pixel = 132;
			13586: Pixel = 128;
			13587: Pixel = 122;
			13588: Pixel = 122;
			13589: Pixel = 129;
			13590: Pixel = 154;
			13591: Pixel = 190;
			13592: Pixel = 225;
			13593: Pixel = 198;
			13594: Pixel = 155;
			13595: Pixel = 154;
			13596: Pixel = 147;
			13597: Pixel = 141;
			13598: Pixel = 133;
			13599: Pixel = 129;
			13600: Pixel = 110;
			13601: Pixel = 61;
			13602: Pixel = 42;
			13603: Pixel = 53;
			13604: Pixel = 65;
			13605: Pixel = 79;
			13606: Pixel = 43;
			13607: Pixel = 46;
			13608: Pixel = 145;
			13609: Pixel = 157;
			13610: Pixel = 121;
			13611: Pixel = 36;
			13612: Pixel = 50;
			13613: Pixel = 41;
			13614: Pixel = 76;
			13615: Pixel = 139;
			13616: Pixel = 137;
			13617: Pixel = 150;
			13618: Pixel = 161;
			13619: Pixel = 158;
			13620: Pixel = 154;
			13621: Pixel = 153;
			13622: Pixel = 154;
			13623: Pixel = 153;
			13624: Pixel = 151;
			13625: Pixel = 150;
			13626: Pixel = 148;
			13627: Pixel = 147;
			13628: Pixel = 147;
			13629: Pixel = 145;
			13630: Pixel = 143;
			13631: Pixel = 140;
			13632: Pixel = 139;
			13633: Pixel = 138;
			13634: Pixel = 130;
			13635: Pixel = 139;
			13636: Pixel = 177;
			13637: Pixel = 194;
			13638: Pixel = 195;
			13639: Pixel = 192;
			13640: Pixel = 192;
			13641: Pixel = 192;
			13642: Pixel = 197;
			13643: Pixel = 203;
			13644: Pixel = 206;
			13645: Pixel = 209;
			13646: Pixel = 209;
			13647: Pixel = 206;
			13648: Pixel = 202;
			13649: Pixel = 202;
			13650: Pixel = 81;
			13651: Pixel = 78;
			13652: Pixel = 73;
			13653: Pixel = 73;
			13654: Pixel = 71;
			13655: Pixel = 61;
			13656: Pixel = 51;
			13657: Pixel = 46;
			13658: Pixel = 92;
			13659: Pixel = 136;
			13660: Pixel = 157;
			13661: Pixel = 169;
			13662: Pixel = 173;
			13663: Pixel = 174;
			13664: Pixel = 175;
			13665: Pixel = 176;
			13666: Pixel = 166;
			13667: Pixel = 150;
			13668: Pixel = 118;
			13669: Pixel = 80;
			13670: Pixel = 74;
			13671: Pixel = 84;
			13672: Pixel = 117;
			13673: Pixel = 123;
			13674: Pixel = 112;
			13675: Pixel = 130;
			13676: Pixel = 93;
			13677: Pixel = 70;
			13678: Pixel = 111;
			13679: Pixel = 84;
			13680: Pixel = 89;
			13681: Pixel = 74;
			13682: Pixel = 82;
			13683: Pixel = 100;
			13684: Pixel = 96;
			13685: Pixel = 91;
			13686: Pixel = 122;
			13687: Pixel = 118;
			13688: Pixel = 85;
			13689: Pixel = 44;
			13690: Pixel = 47;
			13691: Pixel = 49;
			13692: Pixel = 43;
			13693: Pixel = 42;
			13694: Pixel = 56;
			13695: Pixel = 83;
			13696: Pixel = 79;
			13697: Pixel = 90;
			13698: Pixel = 116;
			13699: Pixel = 92;
			13700: Pixel = 143;
			13701: Pixel = 85;
			13702: Pixel = 45;
			13703: Pixel = 43;
			13704: Pixel = 23;
			13705: Pixel = 106;
			13706: Pixel = 123;
			13707: Pixel = 157;
			13708: Pixel = 215;
			13709: Pixel = 126;
			13710: Pixel = 27;
			13711: Pixel = 39;
			13712: Pixel = 42;
			13713: Pixel = 81;
			13714: Pixel = 67;
			13715: Pixel = 88;
			13716: Pixel = 109;
			13717: Pixel = 122;
			13718: Pixel = 126;
			13719: Pixel = 131;
			13720: Pixel = 135;
			13721: Pixel = 139;
			13722: Pixel = 145;
			13723: Pixel = 150;
			13724: Pixel = 152;
			13725: Pixel = 156;
			13726: Pixel = 156;
			13727: Pixel = 160;
			13728: Pixel = 164;
			13729: Pixel = 163;
			13730: Pixel = 162;
			13731: Pixel = 158;
			13732: Pixel = 147;
			13733: Pixel = 136;
			13734: Pixel = 126;
			13735: Pixel = 128;
			13736: Pixel = 129;
			13737: Pixel = 122;
			13738: Pixel = 120;
			13739: Pixel = 129;
			13740: Pixel = 149;
			13741: Pixel = 177;
			13742: Pixel = 225;
			13743: Pixel = 207;
			13744: Pixel = 154;
			13745: Pixel = 153;
			13746: Pixel = 149;
			13747: Pixel = 140;
			13748: Pixel = 132;
			13749: Pixel = 126;
			13750: Pixel = 97;
			13751: Pixel = 48;
			13752: Pixel = 44;
			13753: Pixel = 55;
			13754: Pixel = 67;
			13755: Pixel = 75;
			13756: Pixel = 44;
			13757: Pixel = 40;
			13758: Pixel = 135;
			13759: Pixel = 160;
			13760: Pixel = 128;
			13761: Pixel = 46;
			13762: Pixel = 43;
			13763: Pixel = 44;
			13764: Pixel = 98;
			13765: Pixel = 143;
			13766: Pixel = 137;
			13767: Pixel = 155;
			13768: Pixel = 159;
			13769: Pixel = 157;
			13770: Pixel = 152;
			13771: Pixel = 151;
			13772: Pixel = 152;
			13773: Pixel = 152;
			13774: Pixel = 152;
			13775: Pixel = 150;
			13776: Pixel = 147;
			13777: Pixel = 148;
			13778: Pixel = 147;
			13779: Pixel = 145;
			13780: Pixel = 144;
			13781: Pixel = 141;
			13782: Pixel = 139;
			13783: Pixel = 135;
			13784: Pixel = 130;
			13785: Pixel = 160;
			13786: Pixel = 190;
			13787: Pixel = 196;
			13788: Pixel = 194;
			13789: Pixel = 192;
			13790: Pixel = 193;
			13791: Pixel = 196;
			13792: Pixel = 203;
			13793: Pixel = 208;
			13794: Pixel = 207;
			13795: Pixel = 206;
			13796: Pixel = 207;
			13797: Pixel = 206;
			13798: Pixel = 206;
			13799: Pixel = 205;
			13800: Pixel = 81;
			13801: Pixel = 79;
			13802: Pixel = 77;
			13803: Pixel = 76;
			13804: Pixel = 70;
			13805: Pixel = 59;
			13806: Pixel = 49;
			13807: Pixel = 43;
			13808: Pixel = 89;
			13809: Pixel = 134;
			13810: Pixel = 157;
			13811: Pixel = 169;
			13812: Pixel = 174;
			13813: Pixel = 175;
			13814: Pixel = 177;
			13815: Pixel = 178;
			13816: Pixel = 168;
			13817: Pixel = 150;
			13818: Pixel = 120;
			13819: Pixel = 79;
			13820: Pixel = 69;
			13821: Pixel = 92;
			13822: Pixel = 114;
			13823: Pixel = 114;
			13824: Pixel = 115;
			13825: Pixel = 125;
			13826: Pixel = 79;
			13827: Pixel = 77;
			13828: Pixel = 79;
			13829: Pixel = 107;
			13830: Pixel = 83;
			13831: Pixel = 81;
			13832: Pixel = 73;
			13833: Pixel = 105;
			13834: Pixel = 67;
			13835: Pixel = 91;
			13836: Pixel = 111;
			13837: Pixel = 124;
			13838: Pixel = 78;
			13839: Pixel = 58;
			13840: Pixel = 41;
			13841: Pixel = 56;
			13842: Pixel = 54;
			13843: Pixel = 37;
			13844: Pixel = 54;
			13845: Pixel = 81;
			13846: Pixel = 86;
			13847: Pixel = 131;
			13848: Pixel = 125;
			13849: Pixel = 78;
			13850: Pixel = 79;
			13851: Pixel = 41;
			13852: Pixel = 41;
			13853: Pixel = 37;
			13854: Pixel = 95;
			13855: Pixel = 119;
			13856: Pixel = 109;
			13857: Pixel = 169;
			13858: Pixel = 166;
			13859: Pixel = 62;
			13860: Pixel = 31;
			13861: Pixel = 39;
			13862: Pixel = 45;
			13863: Pixel = 89;
			13864: Pixel = 69;
			13865: Pixel = 85;
			13866: Pixel = 107;
			13867: Pixel = 119;
			13868: Pixel = 126;
			13869: Pixel = 129;
			13870: Pixel = 134;
			13871: Pixel = 137;
			13872: Pixel = 144;
			13873: Pixel = 148;
			13874: Pixel = 152;
			13875: Pixel = 151;
			13876: Pixel = 155;
			13877: Pixel = 158;
			13878: Pixel = 160;
			13879: Pixel = 161;
			13880: Pixel = 160;
			13881: Pixel = 152;
			13882: Pixel = 145;
			13883: Pixel = 127;
			13884: Pixel = 115;
			13885: Pixel = 131;
			13886: Pixel = 136;
			13887: Pixel = 131;
			13888: Pixel = 124;
			13889: Pixel = 129;
			13890: Pixel = 146;
			13891: Pixel = 176;
			13892: Pixel = 222;
			13893: Pixel = 215;
			13894: Pixel = 149;
			13895: Pixel = 148;
			13896: Pixel = 148;
			13897: Pixel = 136;
			13898: Pixel = 129;
			13899: Pixel = 124;
			13900: Pixel = 80;
			13901: Pixel = 39;
			13902: Pixel = 47;
			13903: Pixel = 52;
			13904: Pixel = 71;
			13905: Pixel = 72;
			13906: Pixel = 47;
			13907: Pixel = 35;
			13908: Pixel = 118;
			13909: Pixel = 162;
			13910: Pixel = 143;
			13911: Pixel = 65;
			13912: Pixel = 34;
			13913: Pixel = 52;
			13914: Pixel = 121;
			13915: Pixel = 146;
			13916: Pixel = 141;
			13917: Pixel = 158;
			13918: Pixel = 157;
			13919: Pixel = 154;
			13920: Pixel = 153;
			13921: Pixel = 151;
			13922: Pixel = 150;
			13923: Pixel = 148;
			13924: Pixel = 150;
			13925: Pixel = 150;
			13926: Pixel = 150;
			13927: Pixel = 147;
			13928: Pixel = 147;
			13929: Pixel = 147;
			13930: Pixel = 145;
			13931: Pixel = 141;
			13932: Pixel = 137;
			13933: Pixel = 130;
			13934: Pixel = 139;
			13935: Pixel = 179;
			13936: Pixel = 197;
			13937: Pixel = 196;
			13938: Pixel = 194;
			13939: Pixel = 193;
			13940: Pixel = 195;
			13941: Pixel = 202;
			13942: Pixel = 208;
			13943: Pixel = 207;
			13944: Pixel = 206;
			13945: Pixel = 204;
			13946: Pixel = 206;
			13947: Pixel = 207;
			13948: Pixel = 207;
			13949: Pixel = 206;
			13950: Pixel = 86;
			13951: Pixel = 81;
			13952: Pixel = 79;
			13953: Pixel = 75;
			13954: Pixel = 69;
			13955: Pixel = 63;
			13956: Pixel = 50;
			13957: Pixel = 43;
			13958: Pixel = 92;
			13959: Pixel = 135;
			13960: Pixel = 157;
			13961: Pixel = 170;
			13962: Pixel = 173;
			13963: Pixel = 174;
			13964: Pixel = 176;
			13965: Pixel = 178;
			13966: Pixel = 169;
			13967: Pixel = 150;
			13968: Pixel = 120;
			13969: Pixel = 84;
			13970: Pixel = 95;
			13971: Pixel = 125;
			13972: Pixel = 114;
			13973: Pixel = 102;
			13974: Pixel = 115;
			13975: Pixel = 111;
			13976: Pixel = 70;
			13977: Pixel = 75;
			13978: Pixel = 99;
			13979: Pixel = 107;
			13980: Pixel = 77;
			13981: Pixel = 64;
			13982: Pixel = 81;
			13983: Pixel = 100;
			13984: Pixel = 47;
			13985: Pixel = 106;
			13986: Pixel = 94;
			13987: Pixel = 133;
			13988: Pixel = 73;
			13989: Pixel = 84;
			13990: Pixel = 52;
			13991: Pixel = 56;
			13992: Pixel = 52;
			13993: Pixel = 45;
			13994: Pixel = 46;
			13995: Pixel = 90;
			13996: Pixel = 90;
			13997: Pixel = 51;
			13998: Pixel = 109;
			13999: Pixel = 84;
			14000: Pixel = 37;
			14001: Pixel = 40;
			14002: Pixel = 28;
			14003: Pixel = 80;
			14004: Pixel = 173;
			14005: Pixel = 153;
			14006: Pixel = 140;
			14007: Pixel = 169;
			14008: Pixel = 139;
			14009: Pixel = 43;
			14010: Pixel = 38;
			14011: Pixel = 42;
			14012: Pixel = 46;
			14013: Pixel = 95;
			14014: Pixel = 71;
			14015: Pixel = 86;
			14016: Pixel = 111;
			14017: Pixel = 122;
			14018: Pixel = 127;
			14019: Pixel = 129;
			14020: Pixel = 132;
			14021: Pixel = 139;
			14022: Pixel = 143;
			14023: Pixel = 144;
			14024: Pixel = 149;
			14025: Pixel = 151;
			14026: Pixel = 154;
			14027: Pixel = 156;
			14028: Pixel = 157;
			14029: Pixel = 159;
			14030: Pixel = 158;
			14031: Pixel = 151;
			14032: Pixel = 145;
			14033: Pixel = 120;
			14034: Pixel = 116;
			14035: Pixel = 138;
			14036: Pixel = 141;
			14037: Pixel = 145;
			14038: Pixel = 136;
			14039: Pixel = 122;
			14040: Pixel = 139;
			14041: Pixel = 176;
			14042: Pixel = 213;
			14043: Pixel = 206;
			14044: Pixel = 146;
			14045: Pixel = 147;
			14046: Pixel = 143;
			14047: Pixel = 135;
			14048: Pixel = 128;
			14049: Pixel = 113;
			14050: Pixel = 54;
			14051: Pixel = 40;
			14052: Pixel = 48;
			14053: Pixel = 54;
			14054: Pixel = 69;
			14055: Pixel = 69;
			14056: Pixel = 48;
			14057: Pixel = 34;
			14058: Pixel = 101;
			14059: Pixel = 168;
			14060: Pixel = 146;
			14061: Pixel = 77;
			14062: Pixel = 29;
			14063: Pixel = 59;
			14064: Pixel = 138;
			14065: Pixel = 145;
			14066: Pixel = 146;
			14067: Pixel = 159;
			14068: Pixel = 155;
			14069: Pixel = 154;
			14070: Pixel = 153;
			14071: Pixel = 149;
			14072: Pixel = 150;
			14073: Pixel = 149;
			14074: Pixel = 149;
			14075: Pixel = 148;
			14076: Pixel = 149;
			14077: Pixel = 148;
			14078: Pixel = 148;
			14079: Pixel = 145;
			14080: Pixel = 144;
			14081: Pixel = 140;
			14082: Pixel = 135;
			14083: Pixel = 129;
			14084: Pixel = 155;
			14085: Pixel = 189;
			14086: Pixel = 197;
			14087: Pixel = 194;
			14088: Pixel = 193;
			14089: Pixel = 194;
			14090: Pixel = 200;
			14091: Pixel = 205;
			14092: Pixel = 207;
			14093: Pixel = 206;
			14094: Pixel = 205;
			14095: Pixel = 204;
			14096: Pixel = 206;
			14097: Pixel = 208;
			14098: Pixel = 207;
			14099: Pixel = 206;
			14100: Pixel = 83;
			14101: Pixel = 80;
			14102: Pixel = 79;
			14103: Pixel = 77;
			14104: Pixel = 72;
			14105: Pixel = 65;
			14106: Pixel = 56;
			14107: Pixel = 53;
			14108: Pixel = 101;
			14109: Pixel = 137;
			14110: Pixel = 155;
			14111: Pixel = 168;
			14112: Pixel = 172;
			14113: Pixel = 173;
			14114: Pixel = 176;
			14115: Pixel = 178;
			14116: Pixel = 169;
			14117: Pixel = 149;
			14118: Pixel = 124;
			14119: Pixel = 96;
			14120: Pixel = 89;
			14121: Pixel = 90;
			14122: Pixel = 93;
			14123: Pixel = 102;
			14124: Pixel = 117;
			14125: Pixel = 106;
			14126: Pixel = 70;
			14127: Pixel = 78;
			14128: Pixel = 110;
			14129: Pixel = 115;
			14130: Pixel = 67;
			14131: Pixel = 44;
			14132: Pixel = 123;
			14133: Pixel = 82;
			14134: Pixel = 53;
			14135: Pixel = 96;
			14136: Pixel = 93;
			14137: Pixel = 148;
			14138: Pixel = 84;
			14139: Pixel = 106;
			14140: Pixel = 47;
			14141: Pixel = 54;
			14142: Pixel = 70;
			14143: Pixel = 45;
			14144: Pixel = 35;
			14145: Pixel = 54;
			14146: Pixel = 46;
			14147: Pixel = 76;
			14148: Pixel = 109;
			14149: Pixel = 42;
			14150: Pixel = 39;
			14151: Pixel = 41;
			14152: Pixel = 23;
			14153: Pixel = 132;
			14154: Pixel = 186;
			14155: Pixel = 183;
			14156: Pixel = 193;
			14157: Pixel = 146;
			14158: Pixel = 50;
			14159: Pixel = 30;
			14160: Pixel = 42;
			14161: Pixel = 44;
			14162: Pixel = 44;
			14163: Pixel = 96;
			14164: Pixel = 79;
			14165: Pixel = 91;
			14166: Pixel = 109;
			14167: Pixel = 120;
			14168: Pixel = 124;
			14169: Pixel = 128;
			14170: Pixel = 131;
			14171: Pixel = 138;
			14172: Pixel = 141;
			14173: Pixel = 145;
			14174: Pixel = 149;
			14175: Pixel = 151;
			14176: Pixel = 151;
			14177: Pixel = 153;
			14178: Pixel = 156;
			14179: Pixel = 157;
			14180: Pixel = 157;
			14181: Pixel = 153;
			14182: Pixel = 146;
			14183: Pixel = 127;
			14184: Pixel = 124;
			14185: Pixel = 134;
			14186: Pixel = 83;
			14187: Pixel = 85;
			14188: Pixel = 111;
			14189: Pixel = 116;
			14190: Pixel = 125;
			14191: Pixel = 156;
			14192: Pixel = 199;
			14193: Pixel = 177;
			14194: Pixel = 145;
			14195: Pixel = 147;
			14196: Pixel = 143;
			14197: Pixel = 133;
			14198: Pixel = 129;
			14199: Pixel = 84;
			14200: Pixel = 40;
			14201: Pixel = 45;
			14202: Pixel = 51;
			14203: Pixel = 57;
			14204: Pixel = 69;
			14205: Pixel = 65;
			14206: Pixel = 51;
			14207: Pixel = 36;
			14208: Pixel = 83;
			14209: Pixel = 168;
			14210: Pixel = 144;
			14211: Pixel = 84;
			14212: Pixel = 33;
			14213: Pixel = 79;
			14214: Pixel = 147;
			14215: Pixel = 143;
			14216: Pixel = 151;
			14217: Pixel = 159;
			14218: Pixel = 154;
			14219: Pixel = 153;
			14220: Pixel = 151;
			14221: Pixel = 149;
			14222: Pixel = 150;
			14223: Pixel = 150;
			14224: Pixel = 150;
			14225: Pixel = 148;
			14226: Pixel = 145;
			14227: Pixel = 147;
			14228: Pixel = 145;
			14229: Pixel = 144;
			14230: Pixel = 142;
			14231: Pixel = 140;
			14232: Pixel = 134;
			14233: Pixel = 133;
			14234: Pixel = 169;
			14235: Pixel = 193;
			14236: Pixel = 197;
			14237: Pixel = 194;
			14238: Pixel = 194;
			14239: Pixel = 199;
			14240: Pixel = 204;
			14241: Pixel = 205;
			14242: Pixel = 204;
			14243: Pixel = 206;
			14244: Pixel = 207;
			14245: Pixel = 207;
			14246: Pixel = 208;
			14247: Pixel = 209;
			14248: Pixel = 208;
			14249: Pixel = 206;
			14250: Pixel = 80;
			14251: Pixel = 78;
			14252: Pixel = 77;
			14253: Pixel = 77;
			14254: Pixel = 71;
			14255: Pixel = 67;
			14256: Pixel = 64;
			14257: Pixel = 69;
			14258: Pixel = 112;
			14259: Pixel = 144;
			14260: Pixel = 158;
			14261: Pixel = 168;
			14262: Pixel = 173;
			14263: Pixel = 174;
			14264: Pixel = 176;
			14265: Pixel = 178;
			14266: Pixel = 170;
			14267: Pixel = 151;
			14268: Pixel = 125;
			14269: Pixel = 84;
			14270: Pixel = 72;
			14271: Pixel = 87;
			14272: Pixel = 97;
			14273: Pixel = 104;
			14274: Pixel = 114;
			14275: Pixel = 96;
			14276: Pixel = 84;
			14277: Pixel = 83;
			14278: Pixel = 96;
			14279: Pixel = 102;
			14280: Pixel = 44;
			14281: Pixel = 84;
			14282: Pixel = 113;
			14283: Pixel = 74;
			14284: Pixel = 74;
			14285: Pixel = 89;
			14286: Pixel = 100;
			14287: Pixel = 139;
			14288: Pixel = 107;
			14289: Pixel = 105;
			14290: Pixel = 47;
			14291: Pixel = 46;
			14292: Pixel = 68;
			14293: Pixel = 82;
			14294: Pixel = 39;
			14295: Pixel = 34;
			14296: Pixel = 51;
			14297: Pixel = 122;
			14298: Pixel = 80;
			14299: Pixel = 39;
			14300: Pixel = 55;
			14301: Pixel = 41;
			14302: Pixel = 60;
			14303: Pixel = 145;
			14304: Pixel = 168;
			14305: Pixel = 184;
			14306: Pixel = 175;
			14307: Pixel = 50;
			14308: Pixel = 33;
			14309: Pixel = 46;
			14310: Pixel = 44;
			14311: Pixel = 45;
			14312: Pixel = 47;
			14313: Pixel = 102;
			14314: Pixel = 85;
			14315: Pixel = 96;
			14316: Pixel = 111;
			14317: Pixel = 119;
			14318: Pixel = 123;
			14319: Pixel = 128;
			14320: Pixel = 131;
			14321: Pixel = 135;
			14322: Pixel = 142;
			14323: Pixel = 145;
			14324: Pixel = 148;
			14325: Pixel = 149;
			14326: Pixel = 150;
			14327: Pixel = 154;
			14328: Pixel = 155;
			14329: Pixel = 157;
			14330: Pixel = 158;
			14331: Pixel = 155;
			14332: Pixel = 149;
			14333: Pixel = 139;
			14334: Pixel = 122;
			14335: Pixel = 125;
			14336: Pixel = 104;
			14337: Pixel = 109;
			14338: Pixel = 108;
			14339: Pixel = 100;
			14340: Pixel = 113;
			14341: Pixel = 142;
			14342: Pixel = 185;
			14343: Pixel = 167;
			14344: Pixel = 152;
			14345: Pixel = 144;
			14346: Pixel = 138;
			14347: Pixel = 134;
			14348: Pixel = 120;
			14349: Pixel = 56;
			14350: Pixel = 47;
			14351: Pixel = 46;
			14352: Pixel = 51;
			14353: Pixel = 61;
			14354: Pixel = 71;
			14355: Pixel = 67;
			14356: Pixel = 52;
			14357: Pixel = 41;
			14358: Pixel = 64;
			14359: Pixel = 163;
			14360: Pixel = 146;
			14361: Pixel = 96;
			14362: Pixel = 41;
			14363: Pixel = 109;
			14364: Pixel = 150;
			14365: Pixel = 144;
			14366: Pixel = 154;
			14367: Pixel = 157;
			14368: Pixel = 154;
			14369: Pixel = 151;
			14370: Pixel = 150;
			14371: Pixel = 150;
			14372: Pixel = 148;
			14373: Pixel = 150;
			14374: Pixel = 149;
			14375: Pixel = 147;
			14376: Pixel = 147;
			14377: Pixel = 145;
			14378: Pixel = 143;
			14379: Pixel = 144;
			14380: Pixel = 142;
			14381: Pixel = 140;
			14382: Pixel = 131;
			14383: Pixel = 141;
			14384: Pixel = 179;
			14385: Pixel = 196;
			14386: Pixel = 196;
			14387: Pixel = 195;
			14388: Pixel = 197;
			14389: Pixel = 204;
			14390: Pixel = 207;
			14391: Pixel = 207;
			14392: Pixel = 206;
			14393: Pixel = 206;
			14394: Pixel = 209;
			14395: Pixel = 210;
			14396: Pixel = 209;
			14397: Pixel = 209;
			14398: Pixel = 207;
			14399: Pixel = 206;
			14400: Pixel = 79;
			14401: Pixel = 79;
			14402: Pixel = 75;
			14403: Pixel = 76;
			14404: Pixel = 71;
			14405: Pixel = 67;
			14406: Pixel = 73;
			14407: Pixel = 82;
			14408: Pixel = 120;
			14409: Pixel = 147;
			14410: Pixel = 160;
			14411: Pixel = 167;
			14412: Pixel = 170;
			14413: Pixel = 171;
			14414: Pixel = 175;
			14415: Pixel = 180;
			14416: Pixel = 170;
			14417: Pixel = 151;
			14418: Pixel = 124;
			14419: Pixel = 84;
			14420: Pixel = 76;
			14421: Pixel = 89;
			14422: Pixel = 95;
			14423: Pixel = 106;
			14424: Pixel = 119;
			14425: Pixel = 99;
			14426: Pixel = 54;
			14427: Pixel = 80;
			14428: Pixel = 80;
			14429: Pixel = 50;
			14430: Pixel = 62;
			14431: Pixel = 113;
			14432: Pixel = 71;
			14433: Pixel = 84;
			14434: Pixel = 73;
			14435: Pixel = 95;
			14436: Pixel = 98;
			14437: Pixel = 114;
			14438: Pixel = 128;
			14439: Pixel = 126;
			14440: Pixel = 61;
			14441: Pixel = 31;
			14442: Pixel = 62;
			14443: Pixel = 160;
			14444: Pixel = 82;
			14445: Pixel = 19;
			14446: Pixel = 63;
			14447: Pixel = 93;
			14448: Pixel = 43;
			14449: Pixel = 73;
			14450: Pixel = 96;
			14451: Pixel = 123;
			14452: Pixel = 129;
			14453: Pixel = 106;
			14454: Pixel = 125;
			14455: Pixel = 188;
			14456: Pixel = 76;
			14457: Pixel = 28;
			14458: Pixel = 51;
			14459: Pixel = 67;
			14460: Pixel = 49;
			14461: Pixel = 41;
			14462: Pixel = 49;
			14463: Pixel = 109;
			14464: Pixel = 88;
			14465: Pixel = 97;
			14466: Pixel = 115;
			14467: Pixel = 119;
			14468: Pixel = 124;
			14469: Pixel = 127;
			14470: Pixel = 129;
			14471: Pixel = 134;
			14472: Pixel = 138;
			14473: Pixel = 144;
			14474: Pixel = 145;
			14475: Pixel = 146;
			14476: Pixel = 148;
			14477: Pixel = 152;
			14478: Pixel = 153;
			14479: Pixel = 156;
			14480: Pixel = 158;
			14481: Pixel = 156;
			14482: Pixel = 153;
			14483: Pixel = 148;
			14484: Pixel = 139;
			14485: Pixel = 130;
			14486: Pixel = 132;
			14487: Pixel = 138;
			14488: Pixel = 134;
			14489: Pixel = 129;
			14490: Pixel = 163;
			14491: Pixel = 186;
			14492: Pixel = 183;
			14493: Pixel = 162;
			14494: Pixel = 152;
			14495: Pixel = 145;
			14496: Pixel = 135;
			14497: Pixel = 133;
			14498: Pixel = 91;
			14499: Pixel = 42;
			14500: Pixel = 49;
			14501: Pixel = 47;
			14502: Pixel = 53;
			14503: Pixel = 67;
			14504: Pixel = 79;
			14505: Pixel = 69;
			14506: Pixel = 54;
			14507: Pixel = 44;
			14508: Pixel = 51;
			14509: Pixel = 156;
			14510: Pixel = 147;
			14511: Pixel = 102;
			14512: Pixel = 50;
			14513: Pixel = 128;
			14514: Pixel = 149;
			14515: Pixel = 145;
			14516: Pixel = 157;
			14517: Pixel = 156;
			14518: Pixel = 154;
			14519: Pixel = 152;
			14520: Pixel = 151;
			14521: Pixel = 150;
			14522: Pixel = 149;
			14523: Pixel = 148;
			14524: Pixel = 149;
			14525: Pixel = 149;
			14526: Pixel = 146;
			14527: Pixel = 145;
			14528: Pixel = 145;
			14529: Pixel = 142;
			14530: Pixel = 142;
			14531: Pixel = 138;
			14532: Pixel = 131;
			14533: Pixel = 150;
			14534: Pixel = 187;
			14535: Pixel = 196;
			14536: Pixel = 195;
			14537: Pixel = 197;
			14538: Pixel = 201;
			14539: Pixel = 207;
			14540: Pixel = 207;
			14541: Pixel = 207;
			14542: Pixel = 206;
			14543: Pixel = 207;
			14544: Pixel = 210;
			14545: Pixel = 210;
			14546: Pixel = 209;
			14547: Pixel = 208;
			14548: Pixel = 206;
			14549: Pixel = 208;
			14550: Pixel = 80;
			14551: Pixel = 76;
			14552: Pixel = 77;
			14553: Pixel = 79;
			14554: Pixel = 73;
			14555: Pixel = 68;
			14556: Pixel = 70;
			14557: Pixel = 92;
			14558: Pixel = 125;
			14559: Pixel = 150;
			14560: Pixel = 160;
			14561: Pixel = 166;
			14562: Pixel = 168;
			14563: Pixel = 172;
			14564: Pixel = 175;
			14565: Pixel = 179;
			14566: Pixel = 171;
			14567: Pixel = 153;
			14568: Pixel = 126;
			14569: Pixel = 85;
			14570: Pixel = 76;
			14571: Pixel = 89;
			14572: Pixel = 94;
			14573: Pixel = 100;
			14574: Pixel = 125;
			14575: Pixel = 124;
			14576: Pixel = 42;
			14577: Pixel = 74;
			14578: Pixel = 72;
			14579: Pixel = 71;
			14580: Pixel = 116;
			14581: Pixel = 60;
			14582: Pixel = 54;
			14583: Pixel = 75;
			14584: Pixel = 83;
			14585: Pixel = 107;
			14586: Pixel = 111;
			14587: Pixel = 97;
			14588: Pixel = 116;
			14589: Pixel = 139;
			14590: Pixel = 99;
			14591: Pixel = 45;
			14592: Pixel = 60;
			14593: Pixel = 127;
			14594: Pixel = 88;
			14595: Pixel = 45;
			14596: Pixel = 60;
			14597: Pixel = 53;
			14598: Pixel = 105;
			14599: Pixel = 114;
			14600: Pixel = 144;
			14601: Pixel = 174;
			14602: Pixel = 109;
			14603: Pixel = 102;
			14604: Pixel = 178;
			14605: Pixel = 139;
			14606: Pixel = 36;
			14607: Pixel = 53;
			14608: Pixel = 51;
			14609: Pixel = 58;
			14610: Pixel = 55;
			14611: Pixel = 47;
			14612: Pixel = 49;
			14613: Pixel = 108;
			14614: Pixel = 92;
			14615: Pixel = 98;
			14616: Pixel = 116;
			14617: Pixel = 122;
			14618: Pixel = 124;
			14619: Pixel = 126;
			14620: Pixel = 129;
			14621: Pixel = 134;
			14622: Pixel = 138;
			14623: Pixel = 142;
			14624: Pixel = 143;
			14625: Pixel = 144;
			14626: Pixel = 147;
			14627: Pixel = 153;
			14628: Pixel = 154;
			14629: Pixel = 156;
			14630: Pixel = 159;
			14631: Pixel = 157;
			14632: Pixel = 155;
			14633: Pixel = 152;
			14634: Pixel = 148;
			14635: Pixel = 144;
			14636: Pixel = 137;
			14637: Pixel = 152;
			14638: Pixel = 174;
			14639: Pixel = 158;
			14640: Pixel = 194;
			14641: Pixel = 199;
			14642: Pixel = 183;
			14643: Pixel = 160;
			14644: Pixel = 148;
			14645: Pixel = 142;
			14646: Pixel = 134;
			14647: Pixel = 126;
			14648: Pixel = 63;
			14649: Pixel = 47;
			14650: Pixel = 47;
			14651: Pixel = 48;
			14652: Pixel = 57;
			14653: Pixel = 73;
			14654: Pixel = 80;
			14655: Pixel = 69;
			14656: Pixel = 60;
			14657: Pixel = 52;
			14658: Pixel = 42;
			14659: Pixel = 144;
			14660: Pixel = 149;
			14661: Pixel = 97;
			14662: Pixel = 76;
			14663: Pixel = 139;
			14664: Pixel = 146;
			14665: Pixel = 148;
			14666: Pixel = 157;
			14667: Pixel = 154;
			14668: Pixel = 154;
			14669: Pixel = 151;
			14670: Pixel = 151;
			14671: Pixel = 150;
			14672: Pixel = 148;
			14673: Pixel = 148;
			14674: Pixel = 148;
			14675: Pixel = 147;
			14676: Pixel = 146;
			14677: Pixel = 146;
			14678: Pixel = 145;
			14679: Pixel = 142;
			14680: Pixel = 140;
			14681: Pixel = 134;
			14682: Pixel = 131;
			14683: Pixel = 159;
			14684: Pixel = 191;
			14685: Pixel = 195;
			14686: Pixel = 194;
			14687: Pixel = 199;
			14688: Pixel = 205;
			14689: Pixel = 208;
			14690: Pixel = 207;
			14691: Pixel = 205;
			14692: Pixel = 206;
			14693: Pixel = 208;
			14694: Pixel = 209;
			14695: Pixel = 209;
			14696: Pixel = 210;
			14697: Pixel = 208;
			14698: Pixel = 210;
			14699: Pixel = 210;
			14700: Pixel = 76;
			14701: Pixel = 72;
			14702: Pixel = 75;
			14703: Pixel = 76;
			14704: Pixel = 72;
			14705: Pixel = 61;
			14706: Pixel = 65;
			14707: Pixel = 95;
			14708: Pixel = 129;
			14709: Pixel = 150;
			14710: Pixel = 161;
			14711: Pixel = 167;
			14712: Pixel = 169;
			14713: Pixel = 171;
			14714: Pixel = 177;
			14715: Pixel = 180;
			14716: Pixel = 171;
			14717: Pixel = 153;
			14718: Pixel = 125;
			14719: Pixel = 86;
			14720: Pixel = 74;
			14721: Pixel = 87;
			14722: Pixel = 93;
			14723: Pixel = 110;
			14724: Pixel = 143;
			14725: Pixel = 110;
			14726: Pixel = 59;
			14727: Pixel = 69;
			14728: Pixel = 92;
			14729: Pixel = 115;
			14730: Pixel = 74;
			14731: Pixel = 45;
			14732: Pixel = 55;
			14733: Pixel = 72;
			14734: Pixel = 71;
			14735: Pixel = 83;
			14736: Pixel = 99;
			14737: Pixel = 102;
			14738: Pixel = 97;
			14739: Pixel = 122;
			14740: Pixel = 128;
			14741: Pixel = 71;
			14742: Pixel = 85;
			14743: Pixel = 92;
			14744: Pixel = 67;
			14745: Pixel = 57;
			14746: Pixel = 38;
			14747: Pixel = 96;
			14748: Pixel = 153;
			14749: Pixel = 155;
			14750: Pixel = 188;
			14751: Pixel = 133;
			14752: Pixel = 76;
			14753: Pixel = 133;
			14754: Pixel = 163;
			14755: Pixel = 41;
			14756: Pixel = 46;
			14757: Pixel = 52;
			14758: Pixel = 51;
			14759: Pixel = 59;
			14760: Pixel = 62;
			14761: Pixel = 49;
			14762: Pixel = 47;
			14763: Pixel = 102;
			14764: Pixel = 100;
			14765: Pixel = 100;
			14766: Pixel = 116;
			14767: Pixel = 124;
			14768: Pixel = 126;
			14769: Pixel = 128;
			14770: Pixel = 130;
			14771: Pixel = 136;
			14772: Pixel = 140;
			14773: Pixel = 141;
			14774: Pixel = 139;
			14775: Pixel = 141;
			14776: Pixel = 146;
			14777: Pixel = 151;
			14778: Pixel = 152;
			14779: Pixel = 153;
			14780: Pixel = 155;
			14781: Pixel = 156;
			14782: Pixel = 151;
			14783: Pixel = 150;
			14784: Pixel = 148;
			14785: Pixel = 146;
			14786: Pixel = 147;
			14787: Pixel = 172;
			14788: Pixel = 201;
			14789: Pixel = 174;
			14790: Pixel = 191;
			14791: Pixel = 199;
			14792: Pixel = 184;
			14793: Pixel = 157;
			14794: Pixel = 145;
			14795: Pixel = 141;
			14796: Pixel = 139;
			14797: Pixel = 98;
			14798: Pixel = 45;
			14799: Pixel = 50;
			14800: Pixel = 47;
			14801: Pixel = 49;
			14802: Pixel = 63;
			14803: Pixel = 74;
			14804: Pixel = 76;
			14805: Pixel = 68;
			14806: Pixel = 62;
			14807: Pixel = 50;
			14808: Pixel = 35;
			14809: Pixel = 126;
			14810: Pixel = 158;
			14811: Pixel = 101;
			14812: Pixel = 102;
			14813: Pixel = 145;
			14814: Pixel = 143;
			14815: Pixel = 150;
			14816: Pixel = 157;
			14817: Pixel = 154;
			14818: Pixel = 153;
			14819: Pixel = 150;
			14820: Pixel = 150;
			14821: Pixel = 149;
			14822: Pixel = 148;
			14823: Pixel = 148;
			14824: Pixel = 145;
			14825: Pixel = 144;
			14826: Pixel = 146;
			14827: Pixel = 146;
			14828: Pixel = 145;
			14829: Pixel = 141;
			14830: Pixel = 142;
			14831: Pixel = 135;
			14832: Pixel = 133;
			14833: Pixel = 166;
			14834: Pixel = 193;
			14835: Pixel = 195;
			14836: Pixel = 197;
			14837: Pixel = 203;
			14838: Pixel = 208;
			14839: Pixel = 208;
			14840: Pixel = 206;
			14841: Pixel = 205;
			14842: Pixel = 206;
			14843: Pixel = 208;
			14844: Pixel = 208;
			14845: Pixel = 209;
			14846: Pixel = 210;
			14847: Pixel = 210;
			14848: Pixel = 211;
			14849: Pixel = 211;
			14850: Pixel = 73;
			14851: Pixel = 72;
			14852: Pixel = 70;
			14853: Pixel = 71;
			14854: Pixel = 69;
			14855: Pixel = 62;
			14856: Pixel = 69;
			14857: Pixel = 93;
			14858: Pixel = 128;
			14859: Pixel = 149;
			14860: Pixel = 161;
			14861: Pixel = 168;
			14862: Pixel = 169;
			14863: Pixel = 171;
			14864: Pixel = 176;
			14865: Pixel = 179;
			14866: Pixel = 172;
			14867: Pixel = 154;
			14868: Pixel = 125;
			14869: Pixel = 85;
			14870: Pixel = 73;
			14871: Pixel = 83;
			14872: Pixel = 94;
			14873: Pixel = 133;
			14874: Pixel = 122;
			14875: Pixel = 100;
			14876: Pixel = 59;
			14877: Pixel = 87;
			14878: Pixel = 125;
			14879: Pixel = 57;
			14880: Pixel = 56;
			14881: Pixel = 67;
			14882: Pixel = 59;
			14883: Pixel = 67;
			14884: Pixel = 72;
			14885: Pixel = 69;
			14886: Pixel = 88;
			14887: Pixel = 87;
			14888: Pixel = 82;
			14889: Pixel = 130;
			14890: Pixel = 127;
			14891: Pixel = 88;
			14892: Pixel = 118;
			14893: Pixel = 65;
			14894: Pixel = 46;
			14895: Pixel = 49;
			14896: Pixel = 80;
			14897: Pixel = 125;
			14898: Pixel = 150;
			14899: Pixel = 182;
			14900: Pixel = 174;
			14901: Pixel = 92;
			14902: Pixel = 95;
			14903: Pixel = 154;
			14904: Pixel = 60;
			14905: Pixel = 36;
			14906: Pixel = 54;
			14907: Pixel = 48;
			14908: Pixel = 46;
			14909: Pixel = 59;
			14910: Pixel = 63;
			14911: Pixel = 48;
			14912: Pixel = 42;
			14913: Pixel = 93;
			14914: Pixel = 103;
			14915: Pixel = 96;
			14916: Pixel = 114;
			14917: Pixel = 121;
			14918: Pixel = 126;
			14919: Pixel = 129;
			14920: Pixel = 129;
			14921: Pixel = 135;
			14922: Pixel = 137;
			14923: Pixel = 141;
			14924: Pixel = 139;
			14925: Pixel = 141;
			14926: Pixel = 140;
			14927: Pixel = 143;
			14928: Pixel = 148;
			14929: Pixel = 149;
			14930: Pixel = 149;
			14931: Pixel = 153;
			14932: Pixel = 150;
			14933: Pixel = 147;
			14934: Pixel = 150;
			14935: Pixel = 151;
			14936: Pixel = 154;
			14937: Pixel = 182;
			14938: Pixel = 210;
			14939: Pixel = 178;
			14940: Pixel = 191;
			14941: Pixel = 204;
			14942: Pixel = 181;
			14943: Pixel = 153;
			14944: Pixel = 143;
			14945: Pixel = 140;
			14946: Pixel = 133;
			14947: Pixel = 63;
			14948: Pixel = 43;
			14949: Pixel = 49;
			14950: Pixel = 47;
			14951: Pixel = 52;
			14952: Pixel = 63;
			14953: Pixel = 77;
			14954: Pixel = 75;
			14955: Pixel = 66;
			14956: Pixel = 61;
			14957: Pixel = 48;
			14958: Pixel = 34;
			14959: Pixel = 116;
			14960: Pixel = 153;
			14961: Pixel = 101;
			14962: Pixel = 119;
			14963: Pixel = 144;
			14964: Pixel = 145;
			14965: Pixel = 153;
			14966: Pixel = 154;
			14967: Pixel = 154;
			14968: Pixel = 152;
			14969: Pixel = 151;
			14970: Pixel = 149;
			14971: Pixel = 148;
			14972: Pixel = 147;
			14973: Pixel = 148;
			14974: Pixel = 145;
			14975: Pixel = 145;
			14976: Pixel = 145;
			14977: Pixel = 144;
			14978: Pixel = 145;
			14979: Pixel = 142;
			14980: Pixel = 139;
			14981: Pixel = 132;
			14982: Pixel = 134;
			14983: Pixel = 172;
			14984: Pixel = 195;
			14985: Pixel = 195;
			14986: Pixel = 200;
			14987: Pixel = 207;
			14988: Pixel = 209;
			14989: Pixel = 207;
			14990: Pixel = 206;
			14991: Pixel = 208;
			14992: Pixel = 207;
			14993: Pixel = 207;
			14994: Pixel = 207;
			14995: Pixel = 211;
			14996: Pixel = 211;
			14997: Pixel = 210;
			14998: Pixel = 210;
			14999: Pixel = 211;
			15000: Pixel = 70;
			15001: Pixel = 67;
			15002: Pixel = 68;
			15003: Pixel = 69;
			15004: Pixel = 67;
			15005: Pixel = 64;
			15006: Pixel = 71;
			15007: Pixel = 88;
			15008: Pixel = 123;
			15009: Pixel = 148;
			15010: Pixel = 160;
			15011: Pixel = 167;
			15012: Pixel = 170;
			15013: Pixel = 173;
			15014: Pixel = 176;
			15015: Pixel = 179;
			15016: Pixel = 173;
			15017: Pixel = 155;
			15018: Pixel = 127;
			15019: Pixel = 83;
			15020: Pixel = 72;
			15021: Pixel = 83;
			15022: Pixel = 125;
			15023: Pixel = 113;
			15024: Pixel = 115;
			15025: Pixel = 98;
			15026: Pixel = 67;
			15027: Pixel = 96;
			15028: Pixel = 99;
			15029: Pixel = 49;
			15030: Pixel = 60;
			15031: Pixel = 72;
			15032: Pixel = 70;
			15033: Pixel = 69;
			15034: Pixel = 81;
			15035: Pixel = 66;
			15036: Pixel = 71;
			15037: Pixel = 92;
			15038: Pixel = 59;
			15039: Pixel = 102;
			15040: Pixel = 126;
			15041: Pixel = 137;
			15042: Pixel = 100;
			15043: Pixel = 27;
			15044: Pixel = 62;
			15045: Pixel = 125;
			15046: Pixel = 115;
			15047: Pixel = 119;
			15048: Pixel = 167;
			15049: Pixel = 187;
			15050: Pixel = 111;
			15051: Pixel = 83;
			15052: Pixel = 147;
			15053: Pixel = 90;
			15054: Pixel = 28;
			15055: Pixel = 67;
			15056: Pixel = 58;
			15057: Pixel = 48;
			15058: Pixel = 50;
			15059: Pixel = 56;
			15060: Pixel = 73;
			15061: Pixel = 52;
			15062: Pixel = 40;
			15063: Pixel = 86;
			15064: Pixel = 102;
			15065: Pixel = 89;
			15066: Pixel = 109;
			15067: Pixel = 120;
			15068: Pixel = 126;
			15069: Pixel = 128;
			15070: Pixel = 130;
			15071: Pixel = 135;
			15072: Pixel = 138;
			15073: Pixel = 141;
			15074: Pixel = 140;
			15075: Pixel = 137;
			15076: Pixel = 138;
			15077: Pixel = 141;
			15078: Pixel = 143;
			15079: Pixel = 145;
			15080: Pixel = 143;
			15081: Pixel = 144;
			15082: Pixel = 145;
			15083: Pixel = 144;
			15084: Pixel = 148;
			15085: Pixel = 155;
			15086: Pixel = 160;
			15087: Pixel = 181;
			15088: Pixel = 204;
			15089: Pixel = 193;
			15090: Pixel = 198;
			15091: Pixel = 197;
			15092: Pixel = 186;
			15093: Pixel = 148;
			15094: Pixel = 136;
			15095: Pixel = 143;
			15096: Pixel = 108;
			15097: Pixel = 42;
			15098: Pixel = 47;
			15099: Pixel = 55;
			15100: Pixel = 47;
			15101: Pixel = 54;
			15102: Pixel = 64;
			15103: Pixel = 78;
			15104: Pixel = 74;
			15105: Pixel = 66;
			15106: Pixel = 62;
			15107: Pixel = 51;
			15108: Pixel = 33;
			15109: Pixel = 106;
			15110: Pixel = 157;
			15111: Pixel = 108;
			15112: Pixel = 126;
			15113: Pixel = 143;
			15114: Pixel = 146;
			15115: Pixel = 154;
			15116: Pixel = 154;
			15117: Pixel = 154;
			15118: Pixel = 152;
			15119: Pixel = 152;
			15120: Pixel = 148;
			15121: Pixel = 148;
			15122: Pixel = 148;
			15123: Pixel = 148;
			15124: Pixel = 146;
			15125: Pixel = 146;
			15126: Pixel = 145;
			15127: Pixel = 144;
			15128: Pixel = 144;
			15129: Pixel = 141;
			15130: Pixel = 137;
			15131: Pixel = 129;
			15132: Pixel = 136;
			15133: Pixel = 176;
			15134: Pixel = 195;
			15135: Pixel = 198;
			15136: Pixel = 204;
			15137: Pixel = 209;
			15138: Pixel = 208;
			15139: Pixel = 207;
			15140: Pixel = 208;
			15141: Pixel = 209;
			15142: Pixel = 206;
			15143: Pixel = 206;
			15144: Pixel = 209;
			15145: Pixel = 212;
			15146: Pixel = 212;
			15147: Pixel = 211;
			15148: Pixel = 211;
			15149: Pixel = 211;
			15150: Pixel = 65;
			15151: Pixel = 59;
			15152: Pixel = 64;
			15153: Pixel = 68;
			15154: Pixel = 67;
			15155: Pixel = 62;
			15156: Pixel = 68;
			15157: Pixel = 86;
			15158: Pixel = 124;
			15159: Pixel = 150;
			15160: Pixel = 162;
			15161: Pixel = 169;
			15162: Pixel = 171;
			15163: Pixel = 173;
			15164: Pixel = 178;
			15165: Pixel = 181;
			15166: Pixel = 173;
			15167: Pixel = 155;
			15168: Pixel = 125;
			15169: Pixel = 85;
			15170: Pixel = 66;
			15171: Pixel = 107;
			15172: Pixel = 122;
			15173: Pixel = 89;
			15174: Pixel = 121;
			15175: Pixel = 95;
			15176: Pixel = 45;
			15177: Pixel = 81;
			15178: Pixel = 99;
			15179: Pixel = 52;
			15180: Pixel = 65;
			15181: Pixel = 60;
			15182: Pixel = 62;
			15183: Pixel = 81;
			15184: Pixel = 96;
			15185: Pixel = 87;
			15186: Pixel = 78;
			15187: Pixel = 75;
			15188: Pixel = 91;
			15189: Pixel = 61;
			15190: Pixel = 94;
			15191: Pixel = 135;
			15192: Pixel = 98;
			15193: Pixel = 46;
			15194: Pixel = 107;
			15195: Pixel = 140;
			15196: Pixel = 187;
			15197: Pixel = 188;
			15198: Pixel = 199;
			15199: Pixel = 127;
			15200: Pixel = 82;
			15201: Pixel = 131;
			15202: Pixel = 127;
			15203: Pixel = 31;
			15204: Pixel = 40;
			15205: Pixel = 81;
			15206: Pixel = 59;
			15207: Pixel = 42;
			15208: Pixel = 52;
			15209: Pixel = 59;
			15210: Pixel = 75;
			15211: Pixel = 54;
			15212: Pixel = 41;
			15213: Pixel = 83;
			15214: Pixel = 97;
			15215: Pixel = 84;
			15216: Pixel = 102;
			15217: Pixel = 118;
			15218: Pixel = 126;
			15219: Pixel = 130;
			15220: Pixel = 128;
			15221: Pixel = 133;
			15222: Pixel = 135;
			15223: Pixel = 137;
			15224: Pixel = 141;
			15225: Pixel = 137;
			15226: Pixel = 138;
			15227: Pixel = 139;
			15228: Pixel = 131;
			15229: Pixel = 134;
			15230: Pixel = 139;
			15231: Pixel = 142;
			15232: Pixel = 143;
			15233: Pixel = 142;
			15234: Pixel = 144;
			15235: Pixel = 147;
			15236: Pixel = 144;
			15237: Pixel = 141;
			15238: Pixel = 150;
			15239: Pixel = 169;
			15240: Pixel = 157;
			15241: Pixel = 145;
			15242: Pixel = 150;
			15243: Pixel = 121;
			15244: Pixel = 132;
			15245: Pixel = 141;
			15246: Pixel = 69;
			15247: Pixel = 41;
			15248: Pixel = 50;
			15249: Pixel = 53;
			15250: Pixel = 49;
			15251: Pixel = 55;
			15252: Pixel = 67;
			15253: Pixel = 75;
			15254: Pixel = 77;
			15255: Pixel = 73;
			15256: Pixel = 66;
			15257: Pixel = 52;
			15258: Pixel = 29;
			15259: Pixel = 93;
			15260: Pixel = 155;
			15261: Pixel = 113;
			15262: Pixel = 135;
			15263: Pixel = 145;
			15264: Pixel = 145;
			15265: Pixel = 155;
			15266: Pixel = 155;
			15267: Pixel = 153;
			15268: Pixel = 150;
			15269: Pixel = 149;
			15270: Pixel = 147;
			15271: Pixel = 146;
			15272: Pixel = 150;
			15273: Pixel = 147;
			15274: Pixel = 148;
			15275: Pixel = 144;
			15276: Pixel = 145;
			15277: Pixel = 144;
			15278: Pixel = 143;
			15279: Pixel = 140;
			15280: Pixel = 138;
			15281: Pixel = 128;
			15282: Pixel = 137;
			15283: Pixel = 178;
			15284: Pixel = 196;
			15285: Pixel = 203;
			15286: Pixel = 208;
			15287: Pixel = 210;
			15288: Pixel = 208;
			15289: Pixel = 208;
			15290: Pixel = 209;
			15291: Pixel = 209;
			15292: Pixel = 208;
			15293: Pixel = 209;
			15294: Pixel = 211;
			15295: Pixel = 212;
			15296: Pixel = 213;
			15297: Pixel = 211;
			15298: Pixel = 212;
			15299: Pixel = 211;
			15300: Pixel = 57;
			15301: Pixel = 57;
			15302: Pixel = 59;
			15303: Pixel = 65;
			15304: Pixel = 65;
			15305: Pixel = 61;
			15306: Pixel = 70;
			15307: Pixel = 88;
			15308: Pixel = 125;
			15309: Pixel = 151;
			15310: Pixel = 162;
			15311: Pixel = 172;
			15312: Pixel = 174;
			15313: Pixel = 177;
			15314: Pixel = 178;
			15315: Pixel = 179;
			15316: Pixel = 173;
			15317: Pixel = 153;
			15318: Pixel = 125;
			15319: Pixel = 76;
			15320: Pixel = 87;
			15321: Pixel = 131;
			15322: Pixel = 86;
			15323: Pixel = 104;
			15324: Pixel = 147;
			15325: Pixel = 84;
			15326: Pixel = 51;
			15327: Pixel = 70;
			15328: Pixel = 65;
			15329: Pixel = 63;
			15330: Pixel = 67;
			15331: Pixel = 66;
			15332: Pixel = 48;
			15333: Pixel = 81;
			15334: Pixel = 121;
			15335: Pixel = 102;
			15336: Pixel = 98;
			15337: Pixel = 75;
			15338: Pixel = 77;
			15339: Pixel = 100;
			15340: Pixel = 94;
			15341: Pixel = 92;
			15342: Pixel = 93;
			15343: Pixel = 116;
			15344: Pixel = 137;
			15345: Pixel = 144;
			15346: Pixel = 199;
			15347: Pixel = 216;
			15348: Pixel = 145;
			15349: Pixel = 88;
			15350: Pixel = 107;
			15351: Pixel = 162;
			15352: Pixel = 50;
			15353: Pixel = 43;
			15354: Pixel = 43;
			15355: Pixel = 59;
			15356: Pixel = 57;
			15357: Pixel = 43;
			15358: Pixel = 49;
			15359: Pixel = 59;
			15360: Pixel = 72;
			15361: Pixel = 60;
			15362: Pixel = 38;
			15363: Pixel = 81;
			15364: Pixel = 91;
			15365: Pixel = 80;
			15366: Pixel = 95;
			15367: Pixel = 115;
			15368: Pixel = 125;
			15369: Pixel = 131;
			15370: Pixel = 126;
			15371: Pixel = 128;
			15372: Pixel = 133;
			15373: Pixel = 136;
			15374: Pixel = 141;
			15375: Pixel = 142;
			15376: Pixel = 145;
			15377: Pixel = 128;
			15378: Pixel = 90;
			15379: Pixel = 94;
			15380: Pixel = 102;
			15381: Pixel = 113;
			15382: Pixel = 115;
			15383: Pixel = 116;
			15384: Pixel = 107;
			15385: Pixel = 101;
			15386: Pixel = 96;
			15387: Pixel = 102;
			15388: Pixel = 117;
			15389: Pixel = 122;
			15390: Pixel = 96;
			15391: Pixel = 99;
			15392: Pixel = 109;
			15393: Pixel = 113;
			15394: Pixel = 148;
			15395: Pixel = 115;
			15396: Pixel = 43;
			15397: Pixel = 46;
			15398: Pixel = 52;
			15399: Pixel = 47;
			15400: Pixel = 49;
			15401: Pixel = 61;
			15402: Pixel = 67;
			15403: Pixel = 71;
			15404: Pixel = 77;
			15405: Pixel = 70;
			15406: Pixel = 55;
			15407: Pixel = 63;
			15408: Pixel = 33;
			15409: Pixel = 80;
			15410: Pixel = 150;
			15411: Pixel = 126;
			15412: Pixel = 143;
			15413: Pixel = 147;
			15414: Pixel = 147;
			15415: Pixel = 155;
			15416: Pixel = 156;
			15417: Pixel = 151;
			15418: Pixel = 152;
			15419: Pixel = 150;
			15420: Pixel = 149;
			15421: Pixel = 147;
			15422: Pixel = 148;
			15423: Pixel = 147;
			15424: Pixel = 147;
			15425: Pixel = 146;
			15426: Pixel = 143;
			15427: Pixel = 143;
			15428: Pixel = 144;
			15429: Pixel = 143;
			15430: Pixel = 136;
			15431: Pixel = 125;
			15432: Pixel = 141;
			15433: Pixel = 182;
			15434: Pixel = 199;
			15435: Pixel = 207;
			15436: Pixel = 211;
			15437: Pixel = 210;
			15438: Pixel = 209;
			15439: Pixel = 209;
			15440: Pixel = 207;
			15441: Pixel = 208;
			15442: Pixel = 209;
			15443: Pixel = 210;
			15444: Pixel = 211;
			15445: Pixel = 212;
			15446: Pixel = 214;
			15447: Pixel = 212;
			15448: Pixel = 213;
			15449: Pixel = 213;
			15450: Pixel = 55;
			15451: Pixel = 56;
			15452: Pixel = 60;
			15453: Pixel = 65;
			15454: Pixel = 63;
			15455: Pixel = 62;
			15456: Pixel = 78;
			15457: Pixel = 95;
			15458: Pixel = 128;
			15459: Pixel = 151;
			15460: Pixel = 163;
			15461: Pixel = 173;
			15462: Pixel = 176;
			15463: Pixel = 177;
			15464: Pixel = 179;
			15465: Pixel = 181;
			15466: Pixel = 170;
			15467: Pixel = 152;
			15468: Pixel = 119;
			15469: Pixel = 95;
			15470: Pixel = 135;
			15471: Pixel = 94;
			15472: Pixel = 82;
			15473: Pixel = 134;
			15474: Pixel = 138;
			15475: Pixel = 75;
			15476: Pixel = 66;
			15477: Pixel = 56;
			15478: Pixel = 44;
			15479: Pixel = 61;
			15480: Pixel = 66;
			15481: Pixel = 68;
			15482: Pixel = 62;
			15483: Pixel = 82;
			15484: Pixel = 139;
			15485: Pixel = 96;
			15486: Pixel = 99;
			15487: Pixel = 103;
			15488: Pixel = 86;
			15489: Pixel = 103;
			15490: Pixel = 112;
			15491: Pixel = 67;
			15492: Pixel = 69;
			15493: Pixel = 124;
			15494: Pixel = 133;
			15495: Pixel = 147;
			15496: Pixel = 219;
			15497: Pixel = 191;
			15498: Pixel = 98;
			15499: Pixel = 93;
			15500: Pixel = 169;
			15501: Pixel = 94;
			15502: Pixel = 37;
			15503: Pixel = 54;
			15504: Pixel = 43;
			15505: Pixel = 51;
			15506: Pixel = 60;
			15507: Pixel = 44;
			15508: Pixel = 55;
			15509: Pixel = 57;
			15510: Pixel = 65;
			15511: Pixel = 66;
			15512: Pixel = 40;
			15513: Pixel = 76;
			15514: Pixel = 84;
			15515: Pixel = 81;
			15516: Pixel = 90;
			15517: Pixel = 112;
			15518: Pixel = 121;
			15519: Pixel = 126;
			15520: Pixel = 124;
			15521: Pixel = 127;
			15522: Pixel = 132;
			15523: Pixel = 136;
			15524: Pixel = 137;
			15525: Pixel = 146;
			15526: Pixel = 146;
			15527: Pixel = 134;
			15528: Pixel = 123;
			15529: Pixel = 114;
			15530: Pixel = 104;
			15531: Pixel = 104;
			15532: Pixel = 111;
			15533: Pixel = 121;
			15534: Pixel = 120;
			15535: Pixel = 121;
			15536: Pixel = 121;
			15537: Pixel = 128;
			15538: Pixel = 143;
			15539: Pixel = 151;
			15540: Pixel = 138;
			15541: Pixel = 126;
			15542: Pixel = 137;
			15543: Pixel = 142;
			15544: Pixel = 143;
			15545: Pixel = 67;
			15546: Pixel = 41;
			15547: Pixel = 49;
			15548: Pixel = 52;
			15549: Pixel = 45;
			15550: Pixel = 52;
			15551: Pixel = 65;
			15552: Pixel = 61;
			15553: Pixel = 76;
			15554: Pixel = 76;
			15555: Pixel = 71;
			15556: Pixel = 56;
			15557: Pixel = 74;
			15558: Pixel = 38;
			15559: Pixel = 68;
			15560: Pixel = 148;
			15561: Pixel = 141;
			15562: Pixel = 147;
			15563: Pixel = 147;
			15564: Pixel = 150;
			15565: Pixel = 156;
			15566: Pixel = 154;
			15567: Pixel = 151;
			15568: Pixel = 152;
			15569: Pixel = 151;
			15570: Pixel = 151;
			15571: Pixel = 148;
			15572: Pixel = 147;
			15573: Pixel = 145;
			15574: Pixel = 147;
			15575: Pixel = 147;
			15576: Pixel = 144;
			15577: Pixel = 145;
			15578: Pixel = 144;
			15579: Pixel = 141;
			15580: Pixel = 135;
			15581: Pixel = 125;
			15582: Pixel = 146;
			15583: Pixel = 187;
			15584: Pixel = 203;
			15585: Pixel = 210;
			15586: Pixel = 211;
			15587: Pixel = 210;
			15588: Pixel = 210;
			15589: Pixel = 209;
			15590: Pixel = 208;
			15591: Pixel = 210;
			15592: Pixel = 210;
			15593: Pixel = 210;
			15594: Pixel = 211;
			15595: Pixel = 213;
			15596: Pixel = 214;
			15597: Pixel = 212;
			15598: Pixel = 212;
			15599: Pixel = 212;
			15600: Pixel = 55;
			15601: Pixel = 57;
			15602: Pixel = 59;
			15603: Pixel = 63;
			15604: Pixel = 62;
			15605: Pixel = 61;
			15606: Pixel = 82;
			15607: Pixel = 96;
			15608: Pixel = 126;
			15609: Pixel = 150;
			15610: Pixel = 161;
			15611: Pixel = 172;
			15612: Pixel = 176;
			15613: Pixel = 177;
			15614: Pixel = 181;
			15615: Pixel = 180;
			15616: Pixel = 171;
			15617: Pixel = 153;
			15618: Pixel = 126;
			15619: Pixel = 140;
			15620: Pixel = 96;
			15621: Pixel = 69;
			15622: Pixel = 108;
			15623: Pixel = 135;
			15624: Pixel = 109;
			15625: Pixel = 84;
			15626: Pixel = 66;
			15627: Pixel = 83;
			15628: Pixel = 49;
			15629: Pixel = 39;
			15630: Pixel = 67;
			15631: Pixel = 71;
			15632: Pixel = 66;
			15633: Pixel = 88;
			15634: Pixel = 152;
			15635: Pixel = 66;
			15636: Pixel = 85;
			15637: Pixel = 109;
			15638: Pixel = 101;
			15639: Pixel = 78;
			15640: Pixel = 66;
			15641: Pixel = 97;
			15642: Pixel = 115;
			15643: Pixel = 146;
			15644: Pixel = 140;
			15645: Pixel = 123;
			15646: Pixel = 198;
			15647: Pixel = 127;
			15648: Pixel = 100;
			15649: Pixel = 167;
			15650: Pixel = 135;
			15651: Pixel = 39;
			15652: Pixel = 54;
			15653: Pixel = 52;
			15654: Pixel = 43;
			15655: Pixel = 47;
			15656: Pixel = 56;
			15657: Pixel = 46;
			15658: Pixel = 53;
			15659: Pixel = 59;
			15660: Pixel = 62;
			15661: Pixel = 67;
			15662: Pixel = 46;
			15663: Pixel = 70;
			15664: Pixel = 77;
			15665: Pixel = 77;
			15666: Pixel = 81;
			15667: Pixel = 106;
			15668: Pixel = 115;
			15669: Pixel = 120;
			15670: Pixel = 122;
			15671: Pixel = 124;
			15672: Pixel = 127;
			15673: Pixel = 131;
			15674: Pixel = 136;
			15675: Pixel = 144;
			15676: Pixel = 145;
			15677: Pixel = 148;
			15678: Pixel = 138;
			15679: Pixel = 130;
			15680: Pixel = 128;
			15681: Pixel = 128;
			15682: Pixel = 125;
			15683: Pixel = 130;
			15684: Pixel = 139;
			15685: Pixel = 161;
			15686: Pixel = 177;
			15687: Pixel = 178;
			15688: Pixel = 185;
			15689: Pixel = 195;
			15690: Pixel = 155;
			15691: Pixel = 136;
			15692: Pixel = 147;
			15693: Pixel = 148;
			15694: Pixel = 99;
			15695: Pixel = 39;
			15696: Pixel = 46;
			15697: Pixel = 51;
			15698: Pixel = 48;
			15699: Pixel = 42;
			15700: Pixel = 55;
			15701: Pixel = 53;
			15702: Pixel = 61;
			15703: Pixel = 81;
			15704: Pixel = 77;
			15705: Pixel = 69;
			15706: Pixel = 61;
			15707: Pixel = 76;
			15708: Pixel = 41;
			15709: Pixel = 63;
			15710: Pixel = 149;
			15711: Pixel = 147;
			15712: Pixel = 149;
			15713: Pixel = 148;
			15714: Pixel = 151;
			15715: Pixel = 156;
			15716: Pixel = 154;
			15717: Pixel = 153;
			15718: Pixel = 152;
			15719: Pixel = 152;
			15720: Pixel = 152;
			15721: Pixel = 150;
			15722: Pixel = 149;
			15723: Pixel = 147;
			15724: Pixel = 147;
			15725: Pixel = 145;
			15726: Pixel = 145;
			15727: Pixel = 145;
			15728: Pixel = 144;
			15729: Pixel = 141;
			15730: Pixel = 134;
			15731: Pixel = 124;
			15732: Pixel = 149;
			15733: Pixel = 193;
			15734: Pixel = 209;
			15735: Pixel = 212;
			15736: Pixel = 211;
			15737: Pixel = 210;
			15738: Pixel = 210;
			15739: Pixel = 210;
			15740: Pixel = 210;
			15741: Pixel = 211;
			15742: Pixel = 212;
			15743: Pixel = 213;
			15744: Pixel = 213;
			15745: Pixel = 213;
			15746: Pixel = 211;
			15747: Pixel = 210;
			15748: Pixel = 210;
			15749: Pixel = 209;
			15750: Pixel = 55;
			15751: Pixel = 54;
			15752: Pixel = 57;
			15753: Pixel = 59;
			15754: Pixel = 58;
			15755: Pixel = 58;
			15756: Pixel = 81;
			15757: Pixel = 94;
			15758: Pixel = 123;
			15759: Pixel = 150;
			15760: Pixel = 161;
			15761: Pixel = 170;
			15762: Pixel = 177;
			15763: Pixel = 178;
			15764: Pixel = 180;
			15765: Pixel = 180;
			15766: Pixel = 171;
			15767: Pixel = 166;
			15768: Pixel = 144;
			15769: Pixel = 92;
			15770: Pixel = 62;
			15771: Pixel = 83;
			15772: Pixel = 136;
			15773: Pixel = 115;
			15774: Pixel = 102;
			15775: Pixel = 64;
			15776: Pixel = 91;
			15777: Pixel = 101;
			15778: Pixel = 41;
			15779: Pixel = 44;
			15780: Pixel = 82;
			15781: Pixel = 76;
			15782: Pixel = 73;
			15783: Pixel = 109;
			15784: Pixel = 147;
			15785: Pixel = 84;
			15786: Pixel = 70;
			15787: Pixel = 83;
			15788: Pixel = 108;
			15789: Pixel = 104;
			15790: Pixel = 84;
			15791: Pixel = 97;
			15792: Pixel = 136;
			15793: Pixel = 153;
			15794: Pixel = 125;
			15795: Pixel = 160;
			15796: Pixel = 162;
			15797: Pixel = 102;
			15798: Pixel = 174;
			15799: Pixel = 149;
			15800: Pixel = 49;
			15801: Pixel = 49;
			15802: Pixel = 52;
			15803: Pixel = 56;
			15804: Pixel = 49;
			15805: Pixel = 46;
			15806: Pixel = 53;
			15807: Pixel = 51;
			15808: Pixel = 49;
			15809: Pixel = 59;
			15810: Pixel = 61;
			15811: Pixel = 69;
			15812: Pixel = 48;
			15813: Pixel = 66;
			15814: Pixel = 79;
			15815: Pixel = 71;
			15816: Pixel = 74;
			15817: Pixel = 100;
			15818: Pixel = 110;
			15819: Pixel = 114;
			15820: Pixel = 117;
			15821: Pixel = 121;
			15822: Pixel = 125;
			15823: Pixel = 128;
			15824: Pixel = 131;
			15825: Pixel = 138;
			15826: Pixel = 142;
			15827: Pixel = 146;
			15828: Pixel = 141;
			15829: Pixel = 134;
			15830: Pixel = 127;
			15831: Pixel = 123;
			15832: Pixel = 126;
			15833: Pixel = 127;
			15834: Pixel = 130;
			15835: Pixel = 143;
			15836: Pixel = 149;
			15837: Pixel = 152;
			15838: Pixel = 145;
			15839: Pixel = 144;
			15840: Pixel = 136;
			15841: Pixel = 145;
			15842: Pixel = 149;
			15843: Pixel = 132;
			15844: Pixel = 57;
			15845: Pixel = 43;
			15846: Pixel = 47;
			15847: Pixel = 52;
			15848: Pixel = 47;
			15849: Pixel = 45;
			15850: Pixel = 57;
			15851: Pixel = 50;
			15852: Pixel = 62;
			15853: Pixel = 82;
			15854: Pixel = 79;
			15855: Pixel = 73;
			15856: Pixel = 63;
			15857: Pixel = 76;
			15858: Pixel = 47;
			15859: Pixel = 63;
			15860: Pixel = 149;
			15861: Pixel = 154;
			15862: Pixel = 152;
			15863: Pixel = 149;
			15864: Pixel = 151;
			15865: Pixel = 156;
			15866: Pixel = 155;
			15867: Pixel = 154;
			15868: Pixel = 153;
			15869: Pixel = 152;
			15870: Pixel = 152;
			15871: Pixel = 151;
			15872: Pixel = 149;
			15873: Pixel = 150;
			15874: Pixel = 147;
			15875: Pixel = 144;
			15876: Pixel = 145;
			15877: Pixel = 144;
			15878: Pixel = 144;
			15879: Pixel = 141;
			15880: Pixel = 133;
			15881: Pixel = 122;
			15882: Pixel = 151;
			15883: Pixel = 199;
			15884: Pixel = 213;
			15885: Pixel = 214;
			15886: Pixel = 212;
			15887: Pixel = 211;
			15888: Pixel = 211;
			15889: Pixel = 213;
			15890: Pixel = 213;
			15891: Pixel = 213;
			15892: Pixel = 214;
			15893: Pixel = 214;
			15894: Pixel = 212;
			15895: Pixel = 209;
			15896: Pixel = 207;
			15897: Pixel = 206;
			15898: Pixel = 205;
			15899: Pixel = 205;
			15900: Pixel = 52;
			15901: Pixel = 50;
			15902: Pixel = 53;
			15903: Pixel = 57;
			15904: Pixel = 54;
			15905: Pixel = 58;
			15906: Pixel = 84;
			15907: Pixel = 90;
			15908: Pixel = 118;
			15909: Pixel = 148;
			15910: Pixel = 159;
			15911: Pixel = 170;
			15912: Pixel = 179;
			15913: Pixel = 178;
			15914: Pixel = 179;
			15915: Pixel = 181;
			15916: Pixel = 172;
			15917: Pixel = 155;
			15918: Pixel = 122;
			15919: Pixel = 76;
			15920: Pixel = 65;
			15921: Pixel = 114;
			15922: Pixel = 130;
			15923: Pixel = 103;
			15924: Pixel = 103;
			15925: Pixel = 46;
			15926: Pixel = 112;
			15927: Pixel = 85;
			15928: Pixel = 38;
			15929: Pixel = 55;
			15930: Pixel = 88;
			15931: Pixel = 60;
			15932: Pixel = 78;
			15933: Pixel = 136;
			15934: Pixel = 117;
			15935: Pixel = 106;
			15936: Pixel = 105;
			15937: Pixel = 95;
			15938: Pixel = 63;
			15939: Pixel = 112;
			15940: Pixel = 129;
			15941: Pixel = 117;
			15942: Pixel = 122;
			15943: Pixel = 154;
			15944: Pixel = 122;
			15945: Pixel = 167;
			15946: Pixel = 158;
			15947: Pixel = 164;
			15948: Pixel = 178;
			15949: Pixel = 63;
			15950: Pixel = 50;
			15951: Pixel = 55;
			15952: Pixel = 55;
			15953: Pixel = 59;
			15954: Pixel = 53;
			15955: Pixel = 53;
			15956: Pixel = 53;
			15957: Pixel = 53;
			15958: Pixel = 59;
			15959: Pixel = 59;
			15960: Pixel = 62;
			15961: Pixel = 69;
			15962: Pixel = 53;
			15963: Pixel = 65;
			15964: Pixel = 78;
			15965: Pixel = 71;
			15966: Pixel = 67;
			15967: Pixel = 86;
			15968: Pixel = 103;
			15969: Pixel = 106;
			15970: Pixel = 112;
			15971: Pixel = 119;
			15972: Pixel = 121;
			15973: Pixel = 128;
			15974: Pixel = 131;
			15975: Pixel = 135;
			15976: Pixel = 137;
			15977: Pixel = 141;
			15978: Pixel = 142;
			15979: Pixel = 136;
			15980: Pixel = 133;
			15981: Pixel = 129;
			15982: Pixel = 127;
			15983: Pixel = 123;
			15984: Pixel = 120;
			15985: Pixel = 123;
			15986: Pixel = 128;
			15987: Pixel = 128;
			15988: Pixel = 124;
			15989: Pixel = 132;
			15990: Pixel = 148;
			15991: Pixel = 147;
			15992: Pixel = 140;
			15993: Pixel = 89;
			15994: Pixel = 45;
			15995: Pixel = 44;
			15996: Pixel = 47;
			15997: Pixel = 49;
			15998: Pixel = 54;
			15999: Pixel = 53;
			16000: Pixel = 56;
			16001: Pixel = 50;
			16002: Pixel = 68;
			16003: Pixel = 79;
			16004: Pixel = 77;
			16005: Pixel = 77;
			16006: Pixel = 61;
			16007: Pixel = 77;
			16008: Pixel = 50;
			16009: Pixel = 59;
			16010: Pixel = 148;
			16011: Pixel = 156;
			16012: Pixel = 152;
			16013: Pixel = 150;
			16014: Pixel = 153;
			16015: Pixel = 154;
			16016: Pixel = 154;
			16017: Pixel = 152;
			16018: Pixel = 153;
			16019: Pixel = 154;
			16020: Pixel = 152;
			16021: Pixel = 151;
			16022: Pixel = 150;
			16023: Pixel = 148;
			16024: Pixel = 148;
			16025: Pixel = 146;
			16026: Pixel = 144;
			16027: Pixel = 142;
			16028: Pixel = 140;
			16029: Pixel = 138;
			16030: Pixel = 131;
			16031: Pixel = 118;
			16032: Pixel = 152;
			16033: Pixel = 203;
			16034: Pixel = 216;
			16035: Pixel = 215;
			16036: Pixel = 212;
			16037: Pixel = 212;
			16038: Pixel = 212;
			16039: Pixel = 215;
			16040: Pixel = 216;
			16041: Pixel = 215;
			16042: Pixel = 213;
			16043: Pixel = 210;
			16044: Pixel = 206;
			16045: Pixel = 205;
			16046: Pixel = 204;
			16047: Pixel = 204;
			16048: Pixel = 205;
			16049: Pixel = 206;
			16050: Pixel = 51;
			16051: Pixel = 51;
			16052: Pixel = 52;
			16053: Pixel = 52;
			16054: Pixel = 48;
			16055: Pixel = 63;
			16056: Pixel = 95;
			16057: Pixel = 91;
			16058: Pixel = 116;
			16059: Pixel = 142;
			16060: Pixel = 154;
			16061: Pixel = 170;
			16062: Pixel = 178;
			16063: Pixel = 178;
			16064: Pixel = 180;
			16065: Pixel = 181;
			16066: Pixel = 171;
			16067: Pixel = 153;
			16068: Pixel = 124;
			16069: Pixel = 79;
			16070: Pixel = 62;
			16071: Pixel = 128;
			16072: Pixel = 108;
			16073: Pixel = 102;
			16074: Pixel = 73;
			16075: Pixel = 48;
			16076: Pixel = 115;
			16077: Pixel = 72;
			16078: Pixel = 37;
			16079: Pixel = 61;
			16080: Pixel = 80;
			16081: Pixel = 45;
			16082: Pixel = 65;
			16083: Pixel = 160;
			16084: Pixel = 123;
			16085: Pixel = 90;
			16086: Pixel = 134;
			16087: Pixel = 111;
			16088: Pixel = 78;
			16089: Pixel = 99;
			16090: Pixel = 131;
			16091: Pixel = 112;
			16092: Pixel = 94;
			16093: Pixel = 120;
			16094: Pixel = 117;
			16095: Pixel = 173;
			16096: Pixel = 172;
			16097: Pixel = 184;
			16098: Pixel = 79;
			16099: Pixel = 42;
			16100: Pixel = 53;
			16101: Pixel = 51;
			16102: Pixel = 55;
			16103: Pixel = 58;
			16104: Pixel = 49;
			16105: Pixel = 50;
			16106: Pixel = 52;
			16107: Pixel = 52;
			16108: Pixel = 58;
			16109: Pixel = 59;
			16110: Pixel = 59;
			16111: Pixel = 61;
			16112: Pixel = 56;
			16113: Pixel = 56;
			16114: Pixel = 70;
			16115: Pixel = 73;
			16116: Pixel = 63;
			16117: Pixel = 79;
			16118: Pixel = 92;
			16119: Pixel = 101;
			16120: Pixel = 105;
			16121: Pixel = 111;
			16122: Pixel = 119;
			16123: Pixel = 125;
			16124: Pixel = 129;
			16125: Pixel = 132;
			16126: Pixel = 136;
			16127: Pixel = 139;
			16128: Pixel = 140;
			16129: Pixel = 137;
			16130: Pixel = 134;
			16131: Pixel = 132;
			16132: Pixel = 131;
			16133: Pixel = 131;
			16134: Pixel = 130;
			16135: Pixel = 124;
			16136: Pixel = 126;
			16137: Pixel = 130;
			16138: Pixel = 139;
			16139: Pixel = 153;
			16140: Pixel = 145;
			16141: Pixel = 145;
			16142: Pixel = 107;
			16143: Pixel = 58;
			16144: Pixel = 48;
			16145: Pixel = 42;
			16146: Pixel = 46;
			16147: Pixel = 51;
			16148: Pixel = 58;
			16149: Pixel = 59;
			16150: Pixel = 53;
			16151: Pixel = 48;
			16152: Pixel = 71;
			16153: Pixel = 84;
			16154: Pixel = 81;
			16155: Pixel = 77;
			16156: Pixel = 60;
			16157: Pixel = 77;
			16158: Pixel = 56;
			16159: Pixel = 56;
			16160: Pixel = 147;
			16161: Pixel = 159;
			16162: Pixel = 152;
			16163: Pixel = 148;
			16164: Pixel = 154;
			16165: Pixel = 154;
			16166: Pixel = 154;
			16167: Pixel = 154;
			16168: Pixel = 153;
			16169: Pixel = 154;
			16170: Pixel = 154;
			16171: Pixel = 156;
			16172: Pixel = 153;
			16173: Pixel = 150;
			16174: Pixel = 149;
			16175: Pixel = 146;
			16176: Pixel = 144;
			16177: Pixel = 142;
			16178: Pixel = 142;
			16179: Pixel = 137;
			16180: Pixel = 128;
			16181: Pixel = 116;
			16182: Pixel = 150;
			16183: Pixel = 206;
			16184: Pixel = 218;
			16185: Pixel = 215;
			16186: Pixel = 213;
			16187: Pixel = 213;
			16188: Pixel = 214;
			16189: Pixel = 215;
			16190: Pixel = 216;
			16191: Pixel = 214;
			16192: Pixel = 209;
			16193: Pixel = 206;
			16194: Pixel = 206;
			16195: Pixel = 207;
			16196: Pixel = 208;
			16197: Pixel = 209;
			16198: Pixel = 210;
			16199: Pixel = 210;
			16200: Pixel = 51;
			16201: Pixel = 51;
			16202: Pixel = 50;
			16203: Pixel = 48;
			16204: Pixel = 44;
			16205: Pixel = 75;
			16206: Pixel = 105;
			16207: Pixel = 101;
			16208: Pixel = 121;
			16209: Pixel = 139;
			16210: Pixel = 151;
			16211: Pixel = 168;
			16212: Pixel = 176;
			16213: Pixel = 177;
			16214: Pixel = 177;
			16215: Pixel = 180;
			16216: Pixel = 171;
			16217: Pixel = 155;
			16218: Pixel = 127;
			16219: Pixel = 81;
			16220: Pixel = 63;
			16221: Pixel = 115;
			16222: Pixel = 113;
			16223: Pixel = 91;
			16224: Pixel = 72;
			16225: Pixel = 71;
			16226: Pixel = 86;
			16227: Pixel = 55;
			16228: Pixel = 39;
			16229: Pixel = 66;
			16230: Pixel = 71;
			16231: Pixel = 55;
			16232: Pixel = 64;
			16233: Pixel = 151;
			16234: Pixel = 126;
			16235: Pixel = 104;
			16236: Pixel = 134;
			16237: Pixel = 120;
			16238: Pixel = 114;
			16239: Pixel = 89;
			16240: Pixel = 104;
			16241: Pixel = 120;
			16242: Pixel = 79;
			16243: Pixel = 118;
			16244: Pixel = 117;
			16245: Pixel = 187;
			16246: Pixel = 208;
			16247: Pixel = 110;
			16248: Pixel = 37;
			16249: Pixel = 53;
			16250: Pixel = 52;
			16251: Pixel = 48;
			16252: Pixel = 54;
			16253: Pixel = 58;
			16254: Pixel = 50;
			16255: Pixel = 51;
			16256: Pixel = 53;
			16257: Pixel = 52;
			16258: Pixel = 50;
			16259: Pixel = 56;
			16260: Pixel = 57;
			16261: Pixel = 60;
			16262: Pixel = 60;
			16263: Pixel = 49;
			16264: Pixel = 60;
			16265: Pixel = 68;
			16266: Pixel = 59;
			16267: Pixel = 69;
			16268: Pixel = 80;
			16269: Pixel = 93;
			16270: Pixel = 103;
			16271: Pixel = 109;
			16272: Pixel = 116;
			16273: Pixel = 126;
			16274: Pixel = 128;
			16275: Pixel = 133;
			16276: Pixel = 136;
			16277: Pixel = 137;
			16278: Pixel = 138;
			16279: Pixel = 138;
			16280: Pixel = 138;
			16281: Pixel = 140;
			16282: Pixel = 140;
			16283: Pixel = 146;
			16284: Pixel = 153;
			16285: Pixel = 160;
			16286: Pixel = 161;
			16287: Pixel = 156;
			16288: Pixel = 157;
			16289: Pixel = 152;
			16290: Pixel = 144;
			16291: Pixel = 141;
			16292: Pixel = 63;
			16293: Pixel = 59;
			16294: Pixel = 46;
			16295: Pixel = 44;
			16296: Pixel = 49;
			16297: Pixel = 55;
			16298: Pixel = 59;
			16299: Pixel = 56;
			16300: Pixel = 51;
			16301: Pixel = 46;
			16302: Pixel = 73;
			16303: Pixel = 87;
			16304: Pixel = 78;
			16305: Pixel = 78;
			16306: Pixel = 67;
			16307: Pixel = 79;
			16308: Pixel = 56;
			16309: Pixel = 52;
			16310: Pixel = 144;
			16311: Pixel = 166;
			16312: Pixel = 150;
			16313: Pixel = 148;
			16314: Pixel = 155;
			16315: Pixel = 156;
			16316: Pixel = 156;
			16317: Pixel = 152;
			16318: Pixel = 153;
			16319: Pixel = 153;
			16320: Pixel = 152;
			16321: Pixel = 152;
			16322: Pixel = 152;
			16323: Pixel = 149;
			16324: Pixel = 148;
			16325: Pixel = 147;
			16326: Pixel = 144;
			16327: Pixel = 142;
			16328: Pixel = 140;
			16329: Pixel = 134;
			16330: Pixel = 126;
			16331: Pixel = 115;
			16332: Pixel = 150;
			16333: Pixel = 209;
			16334: Pixel = 218;
			16335: Pixel = 217;
			16336: Pixel = 215;
			16337: Pixel = 215;
			16338: Pixel = 215;
			16339: Pixel = 214;
			16340: Pixel = 213;
			16341: Pixel = 210;
			16342: Pixel = 209;
			16343: Pixel = 210;
			16344: Pixel = 212;
			16345: Pixel = 210;
			16346: Pixel = 210;
			16347: Pixel = 210;
			16348: Pixel = 209;
			16349: Pixel = 209;
			16350: Pixel = 47;
			16351: Pixel = 47;
			16352: Pixel = 50;
			16353: Pixel = 49;
			16354: Pixel = 49;
			16355: Pixel = 82;
			16356: Pixel = 105;
			16357: Pixel = 101;
			16358: Pixel = 123;
			16359: Pixel = 139;
			16360: Pixel = 152;
			16361: Pixel = 169;
			16362: Pixel = 175;
			16363: Pixel = 175;
			16364: Pixel = 177;
			16365: Pixel = 179;
			16366: Pixel = 170;
			16367: Pixel = 153;
			16368: Pixel = 125;
			16369: Pixel = 84;
			16370: Pixel = 65;
			16371: Pixel = 94;
			16372: Pixel = 114;
			16373: Pixel = 92;
			16374: Pixel = 71;
			16375: Pixel = 92;
			16376: Pixel = 80;
			16377: Pixel = 51;
			16378: Pixel = 37;
			16379: Pixel = 75;
			16380: Pixel = 63;
			16381: Pixel = 51;
			16382: Pixel = 64;
			16383: Pixel = 123;
			16384: Pixel = 100;
			16385: Pixel = 111;
			16386: Pixel = 124;
			16387: Pixel = 127;
			16388: Pixel = 112;
			16389: Pixel = 89;
			16390: Pixel = 82;
			16391: Pixel = 123;
			16392: Pixel = 119;
			16393: Pixel = 100;
			16394: Pixel = 94;
			16395: Pixel = 178;
			16396: Pixel = 144;
			16397: Pixel = 42;
			16398: Pixel = 51;
			16399: Pixel = 51;
			16400: Pixel = 52;
			16401: Pixel = 49;
			16402: Pixel = 56;
			16403: Pixel = 60;
			16404: Pixel = 47;
			16405: Pixel = 52;
			16406: Pixel = 52;
			16407: Pixel = 53;
			16408: Pixel = 46;
			16409: Pixel = 49;
			16410: Pixel = 56;
			16411: Pixel = 57;
			16412: Pixel = 60;
			16413: Pixel = 49;
			16414: Pixel = 58;
			16415: Pixel = 63;
			16416: Pixel = 55;
			16417: Pixel = 66;
			16418: Pixel = 62;
			16419: Pixel = 75;
			16420: Pixel = 94;
			16421: Pixel = 102;
			16422: Pixel = 109;
			16423: Pixel = 121;
			16424: Pixel = 129;
			16425: Pixel = 132;
			16426: Pixel = 135;
			16427: Pixel = 137;
			16428: Pixel = 140;
			16429: Pixel = 142;
			16430: Pixel = 145;
			16431: Pixel = 153;
			16432: Pixel = 154;
			16433: Pixel = 153;
			16434: Pixel = 165;
			16435: Pixel = 170;
			16436: Pixel = 169;
			16437: Pixel = 161;
			16438: Pixel = 158;
			16439: Pixel = 151;
			16440: Pixel = 154;
			16441: Pixel = 114;
			16442: Pixel = 42;
			16443: Pixel = 59;
			16444: Pixel = 43;
			16445: Pixel = 47;
			16446: Pixel = 51;
			16447: Pixel = 59;
			16448: Pixel = 61;
			16449: Pixel = 56;
			16450: Pixel = 56;
			16451: Pixel = 45;
			16452: Pixel = 82;
			16453: Pixel = 89;
			16454: Pixel = 82;
			16455: Pixel = 78;
			16456: Pixel = 71;
			16457: Pixel = 78;
			16458: Pixel = 63;
			16459: Pixel = 53;
			16460: Pixel = 143;
			16461: Pixel = 167;
			16462: Pixel = 149;
			16463: Pixel = 148;
			16464: Pixel = 158;
			16465: Pixel = 156;
			16466: Pixel = 155;
			16467: Pixel = 154;
			16468: Pixel = 153;
			16469: Pixel = 151;
			16470: Pixel = 151;
			16471: Pixel = 151;
			16472: Pixel = 152;
			16473: Pixel = 150;
			16474: Pixel = 149;
			16475: Pixel = 146;
			16476: Pixel = 142;
			16477: Pixel = 141;
			16478: Pixel = 138;
			16479: Pixel = 135;
			16480: Pixel = 126;
			16481: Pixel = 114;
			16482: Pixel = 158;
			16483: Pixel = 214;
			16484: Pixel = 219;
			16485: Pixel = 218;
			16486: Pixel = 215;
			16487: Pixel = 212;
			16488: Pixel = 212;
			16489: Pixel = 211;
			16490: Pixel = 212;
			16491: Pixel = 213;
			16492: Pixel = 212;
			16493: Pixel = 212;
			16494: Pixel = 211;
			16495: Pixel = 209;
			16496: Pixel = 207;
			16497: Pixel = 206;
			16498: Pixel = 206;
			16499: Pixel = 204;
			16500: Pixel = 46;
			16501: Pixel = 49;
			16502: Pixel = 48;
			16503: Pixel = 47;
			16504: Pixel = 50;
			16505: Pixel = 82;
			16506: Pixel = 102;
			16507: Pixel = 99;
			16508: Pixel = 122;
			16509: Pixel = 139;
			16510: Pixel = 153;
			16511: Pixel = 170;
			16512: Pixel = 176;
			16513: Pixel = 175;
			16514: Pixel = 176;
			16515: Pixel = 178;
			16516: Pixel = 171;
			16517: Pixel = 154;
			16518: Pixel = 125;
			16519: Pixel = 81;
			16520: Pixel = 68;
			16521: Pixel = 91;
			16522: Pixel = 104;
			16523: Pixel = 82;
			16524: Pixel = 61;
			16525: Pixel = 78;
			16526: Pixel = 86;
			16527: Pixel = 53;
			16528: Pixel = 44;
			16529: Pixel = 71;
			16530: Pixel = 63;
			16531: Pixel = 48;
			16532: Pixel = 75;
			16533: Pixel = 120;
			16534: Pixel = 84;
			16535: Pixel = 62;
			16536: Pixel = 96;
			16537: Pixel = 132;
			16538: Pixel = 131;
			16539: Pixel = 119;
			16540: Pixel = 92;
			16541: Pixel = 124;
			16542: Pixel = 131;
			16543: Pixel = 113;
			16544: Pixel = 82;
			16545: Pixel = 129;
			16546: Pixel = 91;
			16547: Pixel = 58;
			16548: Pixel = 50;
			16549: Pixel = 54;
			16550: Pixel = 51;
			16551: Pixel = 50;
			16552: Pixel = 62;
			16553: Pixel = 60;
			16554: Pixel = 46;
			16555: Pixel = 54;
			16556: Pixel = 52;
			16557: Pixel = 50;
			16558: Pixel = 52;
			16559: Pixel = 47;
			16560: Pixel = 51;
			16561: Pixel = 56;
			16562: Pixel = 56;
			16563: Pixel = 55;
			16564: Pixel = 57;
			16565: Pixel = 60;
			16566: Pixel = 58;
			16567: Pixel = 66;
			16568: Pixel = 63;
			16569: Pixel = 48;
			16570: Pixel = 66;
			16571: Pixel = 87;
			16572: Pixel = 97;
			16573: Pixel = 111;
			16574: Pixel = 124;
			16575: Pixel = 129;
			16576: Pixel = 133;
			16577: Pixel = 136;
			16578: Pixel = 143;
			16579: Pixel = 145;
			16580: Pixel = 149;
			16581: Pixel = 158;
			16582: Pixel = 168;
			16583: Pixel = 164;
			16584: Pixel = 165;
			16585: Pixel = 167;
			16586: Pixel = 165;
			16587: Pixel = 171;
			16588: Pixel = 165;
			16589: Pixel = 148;
			16590: Pixel = 153;
			16591: Pixel = 78;
			16592: Pixel = 47;
			16593: Pixel = 59;
			16594: Pixel = 48;
			16595: Pixel = 50;
			16596: Pixel = 53;
			16597: Pixel = 62;
			16598: Pixel = 55;
			16599: Pixel = 53;
			16600: Pixel = 57;
			16601: Pixel = 46;
			16602: Pixel = 86;
			16603: Pixel = 93;
			16604: Pixel = 84;
			16605: Pixel = 78;
			16606: Pixel = 74;
			16607: Pixel = 71;
			16608: Pixel = 69;
			16609: Pixel = 51;
			16610: Pixel = 144;
			16611: Pixel = 168;
			16612: Pixel = 149;
			16613: Pixel = 148;
			16614: Pixel = 158;
			16615: Pixel = 156;
			16616: Pixel = 154;
			16617: Pixel = 150;
			16618: Pixel = 151;
			16619: Pixel = 150;
			16620: Pixel = 150;
			16621: Pixel = 150;
			16622: Pixel = 151;
			16623: Pixel = 149;
			16624: Pixel = 148;
			16625: Pixel = 144;
			16626: Pixel = 141;
			16627: Pixel = 139;
			16628: Pixel = 137;
			16629: Pixel = 133;
			16630: Pixel = 126;
			16631: Pixel = 114;
			16632: Pixel = 170;
			16633: Pixel = 218;
			16634: Pixel = 220;
			16635: Pixel = 217;
			16636: Pixel = 211;
			16637: Pixel = 210;
			16638: Pixel = 211;
			16639: Pixel = 212;
			16640: Pixel = 214;
			16641: Pixel = 214;
			16642: Pixel = 211;
			16643: Pixel = 208;
			16644: Pixel = 206;
			16645: Pixel = 206;
			16646: Pixel = 205;
			16647: Pixel = 206;
			16648: Pixel = 207;
			16649: Pixel = 205;
			16650: Pixel = 48;
			16651: Pixel = 51;
			16652: Pixel = 48;
			16653: Pixel = 46;
			16654: Pixel = 50;
			16655: Pixel = 73;
			16656: Pixel = 92;
			16657: Pixel = 103;
			16658: Pixel = 126;
			16659: Pixel = 139;
			16660: Pixel = 154;
			16661: Pixel = 170;
			16662: Pixel = 175;
			16663: Pixel = 175;
			16664: Pixel = 177;
			16665: Pixel = 178;
			16666: Pixel = 172;
			16667: Pixel = 156;
			16668: Pixel = 125;
			16669: Pixel = 80;
			16670: Pixel = 66;
			16671: Pixel = 86;
			16672: Pixel = 98;
			16673: Pixel = 53;
			16674: Pixel = 50;
			16675: Pixel = 79;
			16676: Pixel = 92;
			16677: Pixel = 51;
			16678: Pixel = 57;
			16679: Pixel = 65;
			16680: Pixel = 60;
			16681: Pixel = 45;
			16682: Pixel = 61;
			16683: Pixel = 133;
			16684: Pixel = 101;
			16685: Pixel = 51;
			16686: Pixel = 72;
			16687: Pixel = 110;
			16688: Pixel = 117;
			16689: Pixel = 134;
			16690: Pixel = 127;
			16691: Pixel = 119;
			16692: Pixel = 140;
			16693: Pixel = 122;
			16694: Pixel = 87;
			16695: Pixel = 79;
			16696: Pixel = 60;
			16697: Pixel = 60;
			16698: Pixel = 50;
			16699: Pixel = 56;
			16700: Pixel = 50;
			16701: Pixel = 50;
			16702: Pixel = 59;
			16703: Pixel = 63;
			16704: Pixel = 47;
			16705: Pixel = 57;
			16706: Pixel = 54;
			16707: Pixel = 51;
			16708: Pixel = 55;
			16709: Pixel = 47;
			16710: Pixel = 48;
			16711: Pixel = 55;
			16712: Pixel = 57;
			16713: Pixel = 56;
			16714: Pixel = 55;
			16715: Pixel = 59;
			16716: Pixel = 60;
			16717: Pixel = 59;
			16718: Pixel = 72;
			16719: Pixel = 50;
			16720: Pixel = 44;
			16721: Pixel = 60;
			16722: Pixel = 79;
			16723: Pixel = 100;
			16724: Pixel = 117;
			16725: Pixel = 123;
			16726: Pixel = 131;
			16727: Pixel = 135;
			16728: Pixel = 139;
			16729: Pixel = 145;
			16730: Pixel = 148;
			16731: Pixel = 151;
			16732: Pixel = 162;
			16733: Pixel = 166;
			16734: Pixel = 169;
			16735: Pixel = 168;
			16736: Pixel = 167;
			16737: Pixel = 171;
			16738: Pixel = 161;
			16739: Pixel = 149;
			16740: Pixel = 140;
			16741: Pixel = 61;
			16742: Pixel = 50;
			16743: Pixel = 56;
			16744: Pixel = 56;
			16745: Pixel = 54;
			16746: Pixel = 53;
			16747: Pixel = 63;
			16748: Pixel = 57;
			16749: Pixel = 51;
			16750: Pixel = 53;
			16751: Pixel = 49;
			16752: Pixel = 90;
			16753: Pixel = 91;
			16754: Pixel = 83;
			16755: Pixel = 76;
			16756: Pixel = 80;
			16757: Pixel = 73;
			16758: Pixel = 73;
			16759: Pixel = 52;
			16760: Pixel = 142;
			16761: Pixel = 168;
			16762: Pixel = 151;
			16763: Pixel = 147;
			16764: Pixel = 152;
			16765: Pixel = 154;
			16766: Pixel = 152;
			16767: Pixel = 148;
			16768: Pixel = 150;
			16769: Pixel = 150;
			16770: Pixel = 150;
			16771: Pixel = 148;
			16772: Pixel = 149;
			16773: Pixel = 148;
			16774: Pixel = 145;
			16775: Pixel = 142;
			16776: Pixel = 139;
			16777: Pixel = 138;
			16778: Pixel = 137;
			16779: Pixel = 131;
			16780: Pixel = 122;
			16781: Pixel = 119;
			16782: Pixel = 181;
			16783: Pixel = 220;
			16784: Pixel = 221;
			16785: Pixel = 214;
			16786: Pixel = 210;
			16787: Pixel = 211;
			16788: Pixel = 212;
			16789: Pixel = 214;
			16790: Pixel = 214;
			16791: Pixel = 212;
			16792: Pixel = 208;
			16793: Pixel = 206;
			16794: Pixel = 205;
			16795: Pixel = 204;
			16796: Pixel = 201;
			16797: Pixel = 198;
			16798: Pixel = 179;
			16799: Pixel = 146;
			16800: Pixel = 46;
			16801: Pixel = 46;
			16802: Pixel = 47;
			16803: Pixel = 44;
			16804: Pixel = 47;
			16805: Pixel = 59;
			16806: Pixel = 90;
			16807: Pixel = 105;
			16808: Pixel = 125;
			16809: Pixel = 141;
			16810: Pixel = 157;
			16811: Pixel = 169;
			16812: Pixel = 172;
			16813: Pixel = 173;
			16814: Pixel = 177;
			16815: Pixel = 178;
			16816: Pixel = 172;
			16817: Pixel = 155;
			16818: Pixel = 125;
			16819: Pixel = 74;
			16820: Pixel = 53;
			16821: Pixel = 113;
			16822: Pixel = 95;
			16823: Pixel = 57;
			16824: Pixel = 51;
			16825: Pixel = 87;
			16826: Pixel = 74;
			16827: Pixel = 57;
			16828: Pixel = 63;
			16829: Pixel = 67;
			16830: Pixel = 54;
			16831: Pixel = 47;
			16832: Pixel = 46;
			16833: Pixel = 131;
			16834: Pixel = 129;
			16835: Pixel = 67;
			16836: Pixel = 78;
			16837: Pixel = 86;
			16838: Pixel = 113;
			16839: Pixel = 110;
			16840: Pixel = 136;
			16841: Pixel = 120;
			16842: Pixel = 137;
			16843: Pixel = 152;
			16844: Pixel = 110;
			16845: Pixel = 123;
			16846: Pixel = 70;
			16847: Pixel = 43;
			16848: Pixel = 52;
			16849: Pixel = 52;
			16850: Pixel = 52;
			16851: Pixel = 52;
			16852: Pixel = 66;
			16853: Pixel = 69;
			16854: Pixel = 45;
			16855: Pixel = 60;
			16856: Pixel = 55;
			16857: Pixel = 50;
			16858: Pixel = 55;
			16859: Pixel = 51;
			16860: Pixel = 50;
			16861: Pixel = 49;
			16862: Pixel = 55;
			16863: Pixel = 60;
			16864: Pixel = 57;
			16865: Pixel = 62;
			16866: Pixel = 61;
			16867: Pixel = 57;
			16868: Pixel = 74;
			16869: Pixel = 68;
			16870: Pixel = 52;
			16871: Pixel = 48;
			16872: Pixel = 57;
			16873: Pixel = 69;
			16874: Pixel = 76;
			16875: Pixel = 84;
			16876: Pixel = 100;
			16877: Pixel = 111;
			16878: Pixel = 121;
			16879: Pixel = 131;
			16880: Pixel = 139;
			16881: Pixel = 146;
			16882: Pixel = 150;
			16883: Pixel = 157;
			16884: Pixel = 166;
			16885: Pixel = 164;
			16886: Pixel = 154;
			16887: Pixel = 154;
			16888: Pixel = 147;
			16889: Pixel = 140;
			16890: Pixel = 124;
			16891: Pixel = 58;
			16892: Pixel = 51;
			16893: Pixel = 58;
			16894: Pixel = 56;
			16895: Pixel = 57;
			16896: Pixel = 54;
			16897: Pixel = 64;
			16898: Pixel = 59;
			16899: Pixel = 55;
			16900: Pixel = 52;
			16901: Pixel = 55;
			16902: Pixel = 90;
			16903: Pixel = 95;
			16904: Pixel = 84;
			16905: Pixel = 79;
			16906: Pixel = 85;
			16907: Pixel = 80;
			16908: Pixel = 75;
			16909: Pixel = 57;
			16910: Pixel = 145;
			16911: Pixel = 163;
			16912: Pixel = 146;
			16913: Pixel = 130;
			16914: Pixel = 135;
			16915: Pixel = 141;
			16916: Pixel = 142;
			16917: Pixel = 147;
			16918: Pixel = 147;
			16919: Pixel = 149;
			16920: Pixel = 150;
			16921: Pixel = 149;
			16922: Pixel = 149;
			16923: Pixel = 147;
			16924: Pixel = 144;
			16925: Pixel = 142;
			16926: Pixel = 140;
			16927: Pixel = 137;
			16928: Pixel = 135;
			16929: Pixel = 131;
			16930: Pixel = 118;
			16931: Pixel = 127;
			16932: Pixel = 193;
			16933: Pixel = 219;
			16934: Pixel = 219;
			16935: Pixel = 213;
			16936: Pixel = 211;
			16937: Pixel = 212;
			16938: Pixel = 212;
			16939: Pixel = 213;
			16940: Pixel = 212;
			16941: Pixel = 209;
			16942: Pixel = 207;
			16943: Pixel = 204;
			16944: Pixel = 201;
			16945: Pixel = 190;
			16946: Pixel = 157;
			16947: Pixel = 107;
			16948: Pixel = 69;
			16949: Pixel = 47;
			16950: Pixel = 45;
			16951: Pixel = 48;
			16952: Pixel = 45;
			16953: Pixel = 43;
			16954: Pixel = 42;
			16955: Pixel = 55;
			16956: Pixel = 87;
			16957: Pixel = 93;
			16958: Pixel = 112;
			16959: Pixel = 141;
			16960: Pixel = 157;
			16961: Pixel = 168;
			16962: Pixel = 173;
			16963: Pixel = 172;
			16964: Pixel = 175;
			16965: Pixel = 177;
			16966: Pixel = 169;
			16967: Pixel = 152;
			16968: Pixel = 114;
			16969: Pixel = 65;
			16970: Pixel = 141;
			16971: Pixel = 142;
			16972: Pixel = 113;
			16973: Pixel = 86;
			16974: Pixel = 38;
			16975: Pixel = 81;
			16976: Pixel = 61;
			16977: Pixel = 60;
			16978: Pixel = 62;
			16979: Pixel = 58;
			16980: Pixel = 47;
			16981: Pixel = 47;
			16982: Pixel = 40;
			16983: Pixel = 117;
			16984: Pixel = 148;
			16985: Pixel = 105;
			16986: Pixel = 79;
			16987: Pixel = 64;
			16988: Pixel = 124;
			16989: Pixel = 98;
			16990: Pixel = 95;
			16991: Pixel = 112;
			16992: Pixel = 143;
			16993: Pixel = 147;
			16994: Pixel = 120;
			16995: Pixel = 152;
			16996: Pixel = 136;
			16997: Pixel = 52;
			16998: Pixel = 43;
			16999: Pixel = 50;
			17000: Pixel = 50;
			17001: Pixel = 53;
			17002: Pixel = 76;
			17003: Pixel = 69;
			17004: Pixel = 40;
			17005: Pixel = 60;
			17006: Pixel = 55;
			17007: Pixel = 48;
			17008: Pixel = 53;
			17009: Pixel = 50;
			17010: Pixel = 49;
			17011: Pixel = 48;
			17012: Pixel = 51;
			17013: Pixel = 57;
			17014: Pixel = 62;
			17015: Pixel = 61;
			17016: Pixel = 63;
			17017: Pixel = 54;
			17018: Pixel = 63;
			17019: Pixel = 80;
			17020: Pixel = 69;
			17021: Pixel = 70;
			17022: Pixel = 84;
			17023: Pixel = 88;
			17024: Pixel = 97;
			17025: Pixel = 108;
			17026: Pixel = 115;
			17027: Pixel = 117;
			17028: Pixel = 125;
			17029: Pixel = 130;
			17030: Pixel = 137;
			17031: Pixel = 147;
			17032: Pixel = 154;
			17033: Pixel = 155;
			17034: Pixel = 162;
			17035: Pixel = 164;
			17036: Pixel = 160;
			17037: Pixel = 160;
			17038: Pixel = 147;
			17039: Pixel = 146;
			17040: Pixel = 127;
			17041: Pixel = 62;
			17042: Pixel = 44;
			17043: Pixel = 52;
			17044: Pixel = 59;
			17045: Pixel = 58;
			17046: Pixel = 55;
			17047: Pixel = 62;
			17048: Pixel = 59;
			17049: Pixel = 51;
			17050: Pixel = 51;
			17051: Pixel = 56;
			17052: Pixel = 87;
			17053: Pixel = 97;
			17054: Pixel = 88;
			17055: Pixel = 81;
			17056: Pixel = 84;
			17057: Pixel = 79;
			17058: Pixel = 71;
			17059: Pixel = 68;
			17060: Pixel = 151;
			17061: Pixel = 161;
			17062: Pixel = 131;
			17063: Pixel = 114;
			17064: Pixel = 114;
			17065: Pixel = 125;
			17066: Pixel = 129;
			17067: Pixel = 133;
			17068: Pixel = 135;
			17069: Pixel = 139;
			17070: Pixel = 144;
			17071: Pixel = 144;
			17072: Pixel = 149;
			17073: Pixel = 147;
			17074: Pixel = 144;
			17075: Pixel = 142;
			17076: Pixel = 139;
			17077: Pixel = 134;
			17078: Pixel = 132;
			17079: Pixel = 126;
			17080: Pixel = 112;
			17081: Pixel = 141;
			17082: Pixel = 206;
			17083: Pixel = 218;
			17084: Pixel = 214;
			17085: Pixel = 210;
			17086: Pixel = 210;
			17087: Pixel = 210;
			17088: Pixel = 210;
			17089: Pixel = 209;
			17090: Pixel = 208;
			17091: Pixel = 205;
			17092: Pixel = 197;
			17093: Pixel = 185;
			17094: Pixel = 151;
			17095: Pixel = 98;
			17096: Pixel = 56;
			17097: Pixel = 35;
			17098: Pixel = 38;
			17099: Pixel = 47;
			17100: Pixel = 52;
			17101: Pixel = 55;
			17102: Pixel = 49;
			17103: Pixel = 41;
			17104: Pixel = 39;
			17105: Pixel = 53;
			17106: Pixel = 77;
			17107: Pixel = 79;
			17108: Pixel = 106;
			17109: Pixel = 140;
			17110: Pixel = 155;
			17111: Pixel = 168;
			17112: Pixel = 173;
			17113: Pixel = 173;
			17114: Pixel = 172;
			17115: Pixel = 175;
			17116: Pixel = 170;
			17117: Pixel = 145;
			17118: Pixel = 110;
			17119: Pixel = 163;
			17120: Pixel = 163;
			17121: Pixel = 68;
			17122: Pixel = 98;
			17123: Pixel = 76;
			17124: Pixel = 37;
			17125: Pixel = 77;
			17126: Pixel = 72;
			17127: Pixel = 63;
			17128: Pixel = 66;
			17129: Pixel = 57;
			17130: Pixel = 57;
			17131: Pixel = 45;
			17132: Pixel = 47;
			17133: Pixel = 115;
			17134: Pixel = 128;
			17135: Pixel = 131;
			17136: Pixel = 83;
			17137: Pixel = 50;
			17138: Pixel = 73;
			17139: Pixel = 95;
			17140: Pixel = 131;
			17141: Pixel = 113;
			17142: Pixel = 105;
			17143: Pixel = 157;
			17144: Pixel = 102;
			17145: Pixel = 67;
			17146: Pixel = 144;
			17147: Pixel = 157;
			17148: Pixel = 59;
			17149: Pixel = 38;
			17150: Pixel = 49;
			17151: Pixel = 52;
			17152: Pixel = 76;
			17153: Pixel = 68;
			17154: Pixel = 39;
			17155: Pixel = 65;
			17156: Pixel = 51;
			17157: Pixel = 47;
			17158: Pixel = 51;
			17159: Pixel = 52;
			17160: Pixel = 48;
			17161: Pixel = 49;
			17162: Pixel = 49;
			17163: Pixel = 54;
			17164: Pixel = 59;
			17165: Pixel = 56;
			17166: Pixel = 59;
			17167: Pixel = 50;
			17168: Pixel = 52;
			17169: Pixel = 74;
			17170: Pixel = 84;
			17171: Pixel = 102;
			17172: Pixel = 119;
			17173: Pixel = 129;
			17174: Pixel = 133;
			17175: Pixel = 135;
			17176: Pixel = 141;
			17177: Pixel = 139;
			17178: Pixel = 137;
			17179: Pixel = 141;
			17180: Pixel = 143;
			17181: Pixel = 151;
			17182: Pixel = 156;
			17183: Pixel = 155;
			17184: Pixel = 154;
			17185: Pixel = 156;
			17186: Pixel = 160;
			17187: Pixel = 164;
			17188: Pixel = 173;
			17189: Pixel = 187;
			17190: Pixel = 191;
			17191: Pixel = 171;
			17192: Pixel = 129;
			17193: Pixel = 79;
			17194: Pixel = 48;
			17195: Pixel = 49;
			17196: Pixel = 53;
			17197: Pixel = 57;
			17198: Pixel = 54;
			17199: Pixel = 47;
			17200: Pixel = 53;
			17201: Pixel = 56;
			17202: Pixel = 85;
			17203: Pixel = 94;
			17204: Pixel = 86;
			17205: Pixel = 83;
			17206: Pixel = 82;
			17207: Pixel = 83;
			17208: Pixel = 71;
			17209: Pixel = 71;
			17210: Pixel = 153;
			17211: Pixel = 155;
			17212: Pixel = 118;
			17213: Pixel = 112;
			17214: Pixel = 109;
			17215: Pixel = 110;
			17216: Pixel = 115;
			17217: Pixel = 118;
			17218: Pixel = 119;
			17219: Pixel = 121;
			17220: Pixel = 125;
			17221: Pixel = 129;
			17222: Pixel = 137;
			17223: Pixel = 140;
			17224: Pixel = 140;
			17225: Pixel = 140;
			17226: Pixel = 138;
			17227: Pixel = 136;
			17228: Pixel = 129;
			17229: Pixel = 123;
			17230: Pixel = 112;
			17231: Pixel = 158;
			17232: Pixel = 213;
			17233: Pixel = 216;
			17234: Pixel = 209;
			17235: Pixel = 208;
			17236: Pixel = 209;
			17237: Pixel = 209;
			17238: Pixel = 208;
			17239: Pixel = 207;
			17240: Pixel = 205;
			17241: Pixel = 197;
			17242: Pixel = 179;
			17243: Pixel = 148;
			17244: Pixel = 79;
			17245: Pixel = 37;
			17246: Pixel = 39;
			17247: Pixel = 46;
			17248: Pixel = 61;
			17249: Pixel = 71;
			17250: Pixel = 63;
			17251: Pixel = 62;
			17252: Pixel = 54;
			17253: Pixel = 50;
			17254: Pixel = 42;
			17255: Pixel = 49;
			17256: Pixel = 70;
			17257: Pixel = 70;
			17258: Pixel = 100;
			17259: Pixel = 135;
			17260: Pixel = 152;
			17261: Pixel = 167;
			17262: Pixel = 172;
			17263: Pixel = 170;
			17264: Pixel = 172;
			17265: Pixel = 175;
			17266: Pixel = 164;
			17267: Pixel = 149;
			17268: Pixel = 174;
			17269: Pixel = 139;
			17270: Pixel = 64;
			17271: Pixel = 64;
			17272: Pixel = 105;
			17273: Pixel = 47;
			17274: Pixel = 35;
			17275: Pixel = 74;
			17276: Pixel = 79;
			17277: Pixel = 56;
			17278: Pixel = 61;
			17279: Pixel = 60;
			17280: Pixel = 85;
			17281: Pixel = 55;
			17282: Pixel = 51;
			17283: Pixel = 89;
			17284: Pixel = 125;
			17285: Pixel = 120;
			17286: Pixel = 123;
			17287: Pixel = 65;
			17288: Pixel = 77;
			17289: Pixel = 134;
			17290: Pixel = 141;
			17291: Pixel = 85;
			17292: Pixel = 95;
			17293: Pixel = 117;
			17294: Pixel = 121;
			17295: Pixel = 78;
			17296: Pixel = 93;
			17297: Pixel = 157;
			17298: Pixel = 143;
			17299: Pixel = 59;
			17300: Pixel = 44;
			17301: Pixel = 59;
			17302: Pixel = 78;
			17303: Pixel = 65;
			17304: Pixel = 43;
			17305: Pixel = 69;
			17306: Pixel = 56;
			17307: Pixel = 52;
			17308: Pixel = 49;
			17309: Pixel = 53;
			17310: Pixel = 51;
			17311: Pixel = 50;
			17312: Pixel = 53;
			17313: Pixel = 52;
			17314: Pixel = 58;
			17315: Pixel = 59;
			17316: Pixel = 57;
			17317: Pixel = 53;
			17318: Pixel = 52;
			17319: Pixel = 75;
			17320: Pixel = 90;
			17321: Pixel = 112;
			17322: Pixel = 125;
			17323: Pixel = 128;
			17324: Pixel = 124;
			17325: Pixel = 126;
			17326: Pixel = 130;
			17327: Pixel = 132;
			17328: Pixel = 135;
			17329: Pixel = 137;
			17330: Pixel = 141;
			17331: Pixel = 147;
			17332: Pixel = 148;
			17333: Pixel = 145;
			17334: Pixel = 144;
			17335: Pixel = 144;
			17336: Pixel = 147;
			17337: Pixel = 161;
			17338: Pixel = 173;
			17339: Pixel = 186;
			17340: Pixel = 197;
			17341: Pixel = 203;
			17342: Pixel = 209;
			17343: Pixel = 194;
			17344: Pixel = 146;
			17345: Pixel = 88;
			17346: Pixel = 50;
			17347: Pixel = 47;
			17348: Pixel = 54;
			17349: Pixel = 49;
			17350: Pixel = 50;
			17351: Pixel = 62;
			17352: Pixel = 92;
			17353: Pixel = 94;
			17354: Pixel = 82;
			17355: Pixel = 82;
			17356: Pixel = 80;
			17357: Pixel = 84;
			17358: Pixel = 75;
			17359: Pixel = 78;
			17360: Pixel = 158;
			17361: Pixel = 146;
			17362: Pixel = 120;
			17363: Pixel = 125;
			17364: Pixel = 124;
			17365: Pixel = 115;
			17366: Pixel = 115;
			17367: Pixel = 112;
			17368: Pixel = 111;
			17369: Pixel = 109;
			17370: Pixel = 109;
			17371: Pixel = 111;
			17372: Pixel = 114;
			17373: Pixel = 120;
			17374: Pixel = 123;
			17375: Pixel = 125;
			17376: Pixel = 129;
			17377: Pixel = 129;
			17378: Pixel = 127;
			17379: Pixel = 122;
			17380: Pixel = 113;
			17381: Pixel = 166;
			17382: Pixel = 213;
			17383: Pixel = 211;
			17384: Pixel = 205;
			17385: Pixel = 206;
			17386: Pixel = 208;
			17387: Pixel = 209;
			17388: Pixel = 209;
			17389: Pixel = 204;
			17390: Pixel = 194;
			17391: Pixel = 187;
			17392: Pixel = 163;
			17393: Pixel = 95;
			17394: Pixel = 44;
			17395: Pixel = 45;
			17396: Pixel = 52;
			17397: Pixel = 68;
			17398: Pixel = 83;
			17399: Pixel = 80;
			17400: Pixel = 107;
			17401: Pixel = 88;
			17402: Pixel = 69;
			17403: Pixel = 59;
			17404: Pixel = 50;
			17405: Pixel = 58;
			17406: Pixel = 62;
			17407: Pixel = 55;
			17408: Pixel = 79;
			17409: Pixel = 121;
			17410: Pixel = 149;
			17411: Pixel = 167;
			17412: Pixel = 170;
			17413: Pixel = 170;
			17414: Pixel = 170;
			17415: Pixel = 173;
			17416: Pixel = 175;
			17417: Pixel = 178;
			17418: Pixel = 147;
			17419: Pixel = 65;
			17420: Pixel = 68;
			17421: Pixel = 113;
			17422: Pixel = 103;
			17423: Pixel = 33;
			17424: Pixel = 39;
			17425: Pixel = 53;
			17426: Pixel = 77;
			17427: Pixel = 59;
			17428: Pixel = 52;
			17429: Pixel = 52;
			17430: Pixel = 97;
			17431: Pixel = 73;
			17432: Pixel = 64;
			17433: Pixel = 46;
			17434: Pixel = 94;
			17435: Pixel = 126;
			17436: Pixel = 96;
			17437: Pixel = 104;
			17438: Pixel = 120;
			17439: Pixel = 150;
			17440: Pixel = 96;
			17441: Pixel = 80;
			17442: Pixel = 97;
			17443: Pixel = 107;
			17444: Pixel = 112;
			17445: Pixel = 89;
			17446: Pixel = 148;
			17447: Pixel = 129;
			17448: Pixel = 104;
			17449: Pixel = 127;
			17450: Pixel = 41;
			17451: Pixel = 53;
			17452: Pixel = 73;
			17453: Pixel = 60;
			17454: Pixel = 41;
			17455: Pixel = 72;
			17456: Pixel = 56;
			17457: Pixel = 50;
			17458: Pixel = 47;
			17459: Pixel = 50;
			17460: Pixel = 54;
			17461: Pixel = 49;
			17462: Pixel = 50;
			17463: Pixel = 49;
			17464: Pixel = 56;
			17465: Pixel = 61;
			17466: Pixel = 58;
			17467: Pixel = 56;
			17468: Pixel = 50;
			17469: Pixel = 70;
			17470: Pixel = 93;
			17471: Pixel = 115;
			17472: Pixel = 121;
			17473: Pixel = 124;
			17474: Pixel = 125;
			17475: Pixel = 124;
			17476: Pixel = 128;
			17477: Pixel = 135;
			17478: Pixel = 136;
			17479: Pixel = 137;
			17480: Pixel = 139;
			17481: Pixel = 143;
			17482: Pixel = 141;
			17483: Pixel = 140;
			17484: Pixel = 141;
			17485: Pixel = 143;
			17486: Pixel = 150;
			17487: Pixel = 165;
			17488: Pixel = 177;
			17489: Pixel = 187;
			17490: Pixel = 195;
			17491: Pixel = 197;
			17492: Pixel = 198;
			17493: Pixel = 204;
			17494: Pixel = 210;
			17495: Pixel = 201;
			17496: Pixel = 154;
			17497: Pixel = 81;
			17498: Pixel = 40;
			17499: Pixel = 38;
			17500: Pixel = 40;
			17501: Pixel = 57;
			17502: Pixel = 86;
			17503: Pixel = 91;
			17504: Pixel = 79;
			17505: Pixel = 79;
			17506: Pixel = 79;
			17507: Pixel = 79;
			17508: Pixel = 66;
			17509: Pixel = 81;
			17510: Pixel = 161;
			17511: Pixel = 140;
			17512: Pixel = 128;
			17513: Pixel = 135;
			17514: Pixel = 136;
			17515: Pixel = 131;
			17516: Pixel = 125;
			17517: Pixel = 120;
			17518: Pixel = 115;
			17519: Pixel = 109;
			17520: Pixel = 105;
			17521: Pixel = 102;
			17522: Pixel = 100;
			17523: Pixel = 101;
			17524: Pixel = 106;
			17525: Pixel = 106;
			17526: Pixel = 106;
			17527: Pixel = 109;
			17528: Pixel = 111;
			17529: Pixel = 106;
			17530: Pixel = 101;
			17531: Pixel = 163;
			17532: Pixel = 209;
			17533: Pixel = 207;
			17534: Pixel = 202;
			17535: Pixel = 206;
			17536: Pixel = 208;
			17537: Pixel = 208;
			17538: Pixel = 209;
			17539: Pixel = 204;
			17540: Pixel = 189;
			17541: Pixel = 151;
			17542: Pixel = 81;
			17543: Pixel = 44;
			17544: Pixel = 47;
			17545: Pixel = 59;
			17546: Pixel = 68;
			17547: Pixel = 82;
			17548: Pixel = 84;
			17549: Pixel = 86;
			17550: Pixel = 133;
			17551: Pixel = 126;
			17552: Pixel = 103;
			17553: Pixel = 82;
			17554: Pixel = 65;
			17555: Pixel = 69;
			17556: Pixel = 58;
			17557: Pixel = 49;
			17558: Pixel = 68;
			17559: Pixel = 112;
			17560: Pixel = 148;
			17561: Pixel = 165;
			17562: Pixel = 169;
			17563: Pixel = 172;
			17564: Pixel = 170;
			17565: Pixel = 177;
			17566: Pixel = 182;
			17567: Pixel = 158;
			17568: Pixel = 117;
			17569: Pixel = 80;
			17570: Pixel = 120;
			17571: Pixel = 144;
			17572: Pixel = 41;
			17573: Pixel = 40;
			17574: Pixel = 42;
			17575: Pixel = 41;
			17576: Pixel = 60;
			17577: Pixel = 98;
			17578: Pixel = 36;
			17579: Pixel = 37;
			17580: Pixel = 93;
			17581: Pixel = 91;
			17582: Pixel = 86;
			17583: Pixel = 57;
			17584: Pixel = 37;
			17585: Pixel = 112;
			17586: Pixel = 123;
			17587: Pixel = 86;
			17588: Pixel = 96;
			17589: Pixel = 115;
			17590: Pixel = 76;
			17591: Pixel = 110;
			17592: Pixel = 100;
			17593: Pixel = 111;
			17594: Pixel = 119;
			17595: Pixel = 111;
			17596: Pixel = 138;
			17597: Pixel = 134;
			17598: Pixel = 59;
			17599: Pixel = 112;
			17600: Pixel = 92;
			17601: Pixel = 45;
			17602: Pixel = 73;
			17603: Pixel = 57;
			17604: Pixel = 38;
			17605: Pixel = 71;
			17606: Pixel = 53;
			17607: Pixel = 49;
			17608: Pixel = 47;
			17609: Pixel = 47;
			17610: Pixel = 57;
			17611: Pixel = 53;
			17612: Pixel = 47;
			17613: Pixel = 51;
			17614: Pixel = 56;
			17615: Pixel = 59;
			17616: Pixel = 67;
			17617: Pixel = 59;
			17618: Pixel = 49;
			17619: Pixel = 61;
			17620: Pixel = 92;
			17621: Pixel = 111;
			17622: Pixel = 117;
			17623: Pixel = 122;
			17624: Pixel = 123;
			17625: Pixel = 127;
			17626: Pixel = 128;
			17627: Pixel = 132;
			17628: Pixel = 135;
			17629: Pixel = 136;
			17630: Pixel = 139;
			17631: Pixel = 140;
			17632: Pixel = 140;
			17633: Pixel = 139;
			17634: Pixel = 143;
			17635: Pixel = 147;
			17636: Pixel = 156;
			17637: Pixel = 168;
			17638: Pixel = 180;
			17639: Pixel = 189;
			17640: Pixel = 192;
			17641: Pixel = 193;
			17642: Pixel = 198;
			17643: Pixel = 200;
			17644: Pixel = 200;
			17645: Pixel = 204;
			17646: Pixel = 214;
			17647: Pixel = 206;
			17648: Pixel = 134;
			17649: Pixel = 48;
			17650: Pixel = 30;
			17651: Pixel = 57;
			17652: Pixel = 82;
			17653: Pixel = 89;
			17654: Pixel = 75;
			17655: Pixel = 77;
			17656: Pixel = 73;
			17657: Pixel = 75;
			17658: Pixel = 66;
			17659: Pixel = 83;
			17660: Pixel = 159;
			17661: Pixel = 139;
			17662: Pixel = 141;
			17663: Pixel = 140;
			17664: Pixel = 139;
			17665: Pixel = 139;
			17666: Pixel = 133;
			17667: Pixel = 131;
			17668: Pixel = 128;
			17669: Pixel = 123;
			17670: Pixel = 115;
			17671: Pixel = 109;
			17672: Pixel = 104;
			17673: Pixel = 98;
			17674: Pixel = 95;
			17675: Pixel = 94;
			17676: Pixel = 91;
			17677: Pixel = 102;
			17678: Pixel = 113;
			17679: Pixel = 96;
			17680: Pixel = 76;
			17681: Pixel = 149;
			17682: Pixel = 208;
			17683: Pixel = 205;
			17684: Pixel = 203;
			17685: Pixel = 209;
			17686: Pixel = 208;
			17687: Pixel = 206;
			17688: Pixel = 203;
			17689: Pixel = 195;
			17690: Pixel = 162;
			17691: Pixel = 79;
			17692: Pixel = 39;
			17693: Pixel = 64;
			17694: Pixel = 73;
			17695: Pixel = 72;
			17696: Pixel = 78;
			17697: Pixel = 84;
			17698: Pixel = 86;
			17699: Pixel = 87;
			17700: Pixel = 136;
			17701: Pixel = 137;
			17702: Pixel = 131;
			17703: Pixel = 113;
			17704: Pixel = 91;
			17705: Pixel = 84;
			17706: Pixel = 68;
			17707: Pixel = 46;
			17708: Pixel = 67;
			17709: Pixel = 111;
			17710: Pixel = 148;
			17711: Pixel = 165;
			17712: Pixel = 168;
			17713: Pixel = 169;
			17714: Pixel = 171;
			17715: Pixel = 172;
			17716: Pixel = 168;
			17717: Pixel = 155;
			17718: Pixel = 122;
			17719: Pixel = 121;
			17720: Pixel = 142;
			17721: Pixel = 95;
			17722: Pixel = 33;
			17723: Pixel = 45;
			17724: Pixel = 40;
			17725: Pixel = 42;
			17726: Pixel = 88;
			17727: Pixel = 114;
			17728: Pixel = 50;
			17729: Pixel = 51;
			17730: Pixel = 118;
			17731: Pixel = 85;
			17732: Pixel = 88;
			17733: Pixel = 52;
			17734: Pixel = 45;
			17735: Pixel = 87;
			17736: Pixel = 83;
			17737: Pixel = 116;
			17738: Pixel = 122;
			17739: Pixel = 83;
			17740: Pixel = 69;
			17741: Pixel = 97;
			17742: Pixel = 121;
			17743: Pixel = 102;
			17744: Pixel = 138;
			17745: Pixel = 132;
			17746: Pixel = 112;
			17747: Pixel = 122;
			17748: Pixel = 94;
			17749: Pixel = 61;
			17750: Pixel = 134;
			17751: Pixel = 61;
			17752: Pixel = 63;
			17753: Pixel = 53;
			17754: Pixel = 42;
			17755: Pixel = 74;
			17756: Pixel = 58;
			17757: Pixel = 54;
			17758: Pixel = 51;
			17759: Pixel = 47;
			17760: Pixel = 56;
			17761: Pixel = 63;
			17762: Pixel = 54;
			17763: Pixel = 51;
			17764: Pixel = 54;
			17765: Pixel = 59;
			17766: Pixel = 71;
			17767: Pixel = 66;
			17768: Pixel = 52;
			17769: Pixel = 62;
			17770: Pixel = 91;
			17771: Pixel = 109;
			17772: Pixel = 116;
			17773: Pixel = 118;
			17774: Pixel = 125;
			17775: Pixel = 128;
			17776: Pixel = 125;
			17777: Pixel = 131;
			17778: Pixel = 139;
			17779: Pixel = 141;
			17780: Pixel = 141;
			17781: Pixel = 139;
			17782: Pixel = 137;
			17783: Pixel = 141;
			17784: Pixel = 145;
			17785: Pixel = 151;
			17786: Pixel = 160;
			17787: Pixel = 171;
			17788: Pixel = 179;
			17789: Pixel = 187;
			17790: Pixel = 189;
			17791: Pixel = 189;
			17792: Pixel = 194;
			17793: Pixel = 195;
			17794: Pixel = 200;
			17795: Pixel = 202;
			17796: Pixel = 202;
			17797: Pixel = 210;
			17798: Pixel = 219;
			17799: Pixel = 174;
			17800: Pixel = 66;
			17801: Pixel = 41;
			17802: Pixel = 67;
			17803: Pixel = 88;
			17804: Pixel = 70;
			17805: Pixel = 72;
			17806: Pixel = 74;
			17807: Pixel = 76;
			17808: Pixel = 58;
			17809: Pixel = 93;
			17810: Pixel = 160;
			17811: Pixel = 137;
			17812: Pixel = 147;
			17813: Pixel = 146;
			17814: Pixel = 143;
			17815: Pixel = 141;
			17816: Pixel = 138;
			17817: Pixel = 137;
			17818: Pixel = 136;
			17819: Pixel = 134;
			17820: Pixel = 127;
			17821: Pixel = 122;
			17822: Pixel = 118;
			17823: Pixel = 110;
			17824: Pixel = 105;
			17825: Pixel = 96;
			17826: Pixel = 91;
			17827: Pixel = 116;
			17828: Pixel = 128;
			17829: Pixel = 102;
			17830: Pixel = 73;
			17831: Pixel = 153;
			17832: Pixel = 210;
			17833: Pixel = 207;
			17834: Pixel = 207;
			17835: Pixel = 212;
			17836: Pixel = 209;
			17837: Pixel = 207;
			17838: Pixel = 190;
			17839: Pixel = 142;
			17840: Pixel = 71;
			17841: Pixel = 43;
			17842: Pixel = 70;
			17843: Pixel = 81;
			17844: Pixel = 77;
			17845: Pixel = 81;
			17846: Pixel = 88;
			17847: Pixel = 92;
			17848: Pixel = 85;
			17849: Pixel = 84;
			17850: Pixel = 130;
			17851: Pixel = 140;
			17852: Pixel = 148;
			17853: Pixel = 138;
			17854: Pixel = 119;
			17855: Pixel = 99;
			17856: Pixel = 74;
			17857: Pixel = 46;
			17858: Pixel = 61;
			17859: Pixel = 114;
			17860: Pixel = 148;
			17861: Pixel = 167;
			17862: Pixel = 171;
			17863: Pixel = 171;
			17864: Pixel = 172;
			17865: Pixel = 175;
			17866: Pixel = 171;
			17867: Pixel = 145;
			17868: Pixel = 150;
			17869: Pixel = 170;
			17870: Pixel = 96;
			17871: Pixel = 70;
			17872: Pixel = 44;
			17873: Pixel = 42;
			17874: Pixel = 38;
			17875: Pixel = 35;
			17876: Pixel = 73;
			17877: Pixel = 96;
			17878: Pixel = 104;
			17879: Pixel = 116;
			17880: Pixel = 91;
			17881: Pixel = 67;
			17882: Pixel = 70;
			17883: Pixel = 70;
			17884: Pixel = 106;
			17885: Pixel = 73;
			17886: Pixel = 61;
			17887: Pixel = 110;
			17888: Pixel = 72;
			17889: Pixel = 56;
			17890: Pixel = 77;
			17891: Pixel = 85;
			17892: Pixel = 105;
			17893: Pixel = 128;
			17894: Pixel = 139;
			17895: Pixel = 139;
			17896: Pixel = 135;
			17897: Pixel = 50;
			17898: Pixel = 120;
			17899: Pixel = 72;
			17900: Pixel = 94;
			17901: Pixel = 110;
			17902: Pixel = 50;
			17903: Pixel = 52;
			17904: Pixel = 44;
			17905: Pixel = 73;
			17906: Pixel = 60;
			17907: Pixel = 53;
			17908: Pixel = 52;
			17909: Pixel = 48;
			17910: Pixel = 55;
			17911: Pixel = 62;
			17912: Pixel = 55;
			17913: Pixel = 50;
			17914: Pixel = 56;
			17915: Pixel = 63;
			17916: Pixel = 71;
			17917: Pixel = 78;
			17918: Pixel = 50;
			17919: Pixel = 62;
			17920: Pixel = 91;
			17921: Pixel = 111;
			17922: Pixel = 117;
			17923: Pixel = 123;
			17924: Pixel = 127;
			17925: Pixel = 121;
			17926: Pixel = 130;
			17927: Pixel = 136;
			17928: Pixel = 139;
			17929: Pixel = 142;
			17930: Pixel = 141;
			17931: Pixel = 138;
			17932: Pixel = 136;
			17933: Pixel = 141;
			17934: Pixel = 148;
			17935: Pixel = 156;
			17936: Pixel = 161;
			17937: Pixel = 167;
			17938: Pixel = 175;
			17939: Pixel = 184;
			17940: Pixel = 185;
			17941: Pixel = 188;
			17942: Pixel = 190;
			17943: Pixel = 192;
			17944: Pixel = 197;
			17945: Pixel = 201;
			17946: Pixel = 204;
			17947: Pixel = 206;
			17948: Pixel = 207;
			17949: Pixel = 220;
			17950: Pixel = 192;
			17951: Pixel = 75;
			17952: Pixel = 45;
			17953: Pixel = 80;
			17954: Pixel = 62;
			17955: Pixel = 64;
			17956: Pixel = 73;
			17957: Pixel = 74;
			17958: Pixel = 49;
			17959: Pixel = 98;
			17960: Pixel = 159;
			17961: Pixel = 138;
			17962: Pixel = 150;
			17963: Pixel = 147;
			17964: Pixel = 145;
			17965: Pixel = 143;
			17966: Pixel = 142;
			17967: Pixel = 141;
			17968: Pixel = 139;
			17969: Pixel = 135;
			17970: Pixel = 134;
			17971: Pixel = 130;
			17972: Pixel = 125;
			17973: Pixel = 121;
			17974: Pixel = 117;
			17975: Pixel = 111;
			17976: Pixel = 103;
			17977: Pixel = 123;
			17978: Pixel = 134;
			17979: Pixel = 101;
			17980: Pixel = 93;
			17981: Pixel = 177;
			17982: Pixel = 211;
			17983: Pixel = 210;
			17984: Pixel = 211;
			17985: Pixel = 212;
			17986: Pixel = 208;
			17987: Pixel = 205;
			17988: Pixel = 168;
			17989: Pixel = 72;
			17990: Pixel = 38;
			17991: Pixel = 72;
			17992: Pixel = 91;
			17993: Pixel = 82;
			17994: Pixel = 78;
			17995: Pixel = 90;
			17996: Pixel = 98;
			17997: Pixel = 96;
			17998: Pixel = 85;
			17999: Pixel = 86;
			18000: Pixel = 128;
			18001: Pixel = 138;
			18002: Pixel = 151;
			18003: Pixel = 150;
			18004: Pixel = 137;
			18005: Pixel = 119;
			18006: Pixel = 86;
			18007: Pixel = 50;
			18008: Pixel = 61;
			18009: Pixel = 112;
			18010: Pixel = 148;
			18011: Pixel = 168;
			18012: Pixel = 175;
			18013: Pixel = 173;
			18014: Pixel = 172;
			18015: Pixel = 176;
			18016: Pixel = 170;
			18017: Pixel = 143;
			18018: Pixel = 188;
			18019: Pixel = 167;
			18020: Pixel = 102;
			18021: Pixel = 59;
			18022: Pixel = 48;
			18023: Pixel = 50;
			18024: Pixel = 51;
			18025: Pixel = 53;
			18026: Pixel = 69;
			18027: Pixel = 40;
			18028: Pixel = 67;
			18029: Pixel = 73;
			18030: Pixel = 54;
			18031: Pixel = 57;
			18032: Pixel = 67;
			18033: Pixel = 81;
			18034: Pixel = 75;
			18035: Pixel = 32;
			18036: Pixel = 102;
			18037: Pixel = 98;
			18038: Pixel = 45;
			18039: Pixel = 76;
			18040: Pixel = 66;
			18041: Pixel = 97;
			18042: Pixel = 89;
			18043: Pixel = 105;
			18044: Pixel = 134;
			18045: Pixel = 136;
			18046: Pixel = 151;
			18047: Pixel = 84;
			18048: Pixel = 79;
			18049: Pixel = 160;
			18050: Pixel = 79;
			18051: Pixel = 127;
			18052: Pixel = 57;
			18053: Pixel = 45;
			18054: Pixel = 46;
			18055: Pixel = 70;
			18056: Pixel = 60;
			18057: Pixel = 53;
			18058: Pixel = 56;
			18059: Pixel = 53;
			18060: Pixel = 56;
			18061: Pixel = 66;
			18062: Pixel = 54;
			18063: Pixel = 52;
			18064: Pixel = 65;
			18065: Pixel = 67;
			18066: Pixel = 77;
			18067: Pixel = 99;
			18068: Pixel = 56;
			18069: Pixel = 51;
			18070: Pixel = 87;
			18071: Pixel = 116;
			18072: Pixel = 119;
			18073: Pixel = 125;
			18074: Pixel = 114;
			18075: Pixel = 126;
			18076: Pixel = 137;
			18077: Pixel = 138;
			18078: Pixel = 136;
			18079: Pixel = 140;
			18080: Pixel = 140;
			18081: Pixel = 138;
			18082: Pixel = 140;
			18083: Pixel = 145;
			18084: Pixel = 151;
			18085: Pixel = 159;
			18086: Pixel = 162;
			18087: Pixel = 166;
			18088: Pixel = 171;
			18089: Pixel = 177;
			18090: Pixel = 180;
			18091: Pixel = 184;
			18092: Pixel = 188;
			18093: Pixel = 191;
			18094: Pixel = 194;
			18095: Pixel = 197;
			18096: Pixel = 202;
			18097: Pixel = 206;
			18098: Pixel = 209;
			18099: Pixel = 209;
			18100: Pixel = 221;
			18101: Pixel = 194;
			18102: Pixel = 72;
			18103: Pixel = 62;
			18104: Pixel = 58;
			18105: Pixel = 60;
			18106: Pixel = 75;
			18107: Pixel = 75;
			18108: Pixel = 49;
			18109: Pixel = 109;
			18110: Pixel = 157;
			18111: Pixel = 137;
			18112: Pixel = 148;
			18113: Pixel = 148;
			18114: Pixel = 145;
			18115: Pixel = 143;
			18116: Pixel = 144;
			18117: Pixel = 143;
			18118: Pixel = 141;
			18119: Pixel = 138;
			18120: Pixel = 137;
			18121: Pixel = 136;
			18122: Pixel = 129;
			18123: Pixel = 128;
			18124: Pixel = 125;
			18125: Pixel = 120;
			18126: Pixel = 114;
			18127: Pixel = 124;
			18128: Pixel = 131;
			18129: Pixel = 109;
			18130: Pixel = 123;
			18131: Pixel = 195;
			18132: Pixel = 211;
			18133: Pixel = 211;
			18134: Pixel = 212;
			18135: Pixel = 212;
			18136: Pixel = 204;
			18137: Pixel = 190;
			18138: Pixel = 133;
			18139: Pixel = 48;
			18140: Pixel = 61;
			18141: Pixel = 92;
			18142: Pixel = 91;
			18143: Pixel = 87;
			18144: Pixel = 87;
			18145: Pixel = 104;
			18146: Pixel = 106;
			18147: Pixel = 94;
			18148: Pixel = 87;
			18149: Pixel = 94;
			18150: Pixel = 102;
			18151: Pixel = 124;
			18152: Pixel = 144;
			18153: Pixel = 153;
			18154: Pixel = 151;
			18155: Pixel = 144;
			18156: Pixel = 104;
			18157: Pixel = 51;
			18158: Pixel = 61;
			18159: Pixel = 112;
			18160: Pixel = 149;
			18161: Pixel = 168;
			18162: Pixel = 176;
			18163: Pixel = 175;
			18164: Pixel = 175;
			18165: Pixel = 177;
			18166: Pixel = 170;
			18167: Pixel = 147;
			18168: Pixel = 170;
			18169: Pixel = 131;
			18170: Pixel = 112;
			18171: Pixel = 43;
			18172: Pixel = 40;
			18173: Pixel = 50;
			18174: Pixel = 51;
			18175: Pixel = 57;
			18176: Pixel = 70;
			18177: Pixel = 58;
			18178: Pixel = 55;
			18179: Pixel = 49;
			18180: Pixel = 64;
			18181: Pixel = 79;
			18182: Pixel = 53;
			18183: Pixel = 35;
			18184: Pixel = 54;
			18185: Pixel = 56;
			18186: Pixel = 59;
			18187: Pixel = 101;
			18188: Pixel = 60;
			18189: Pixel = 63;
			18190: Pixel = 73;
			18191: Pixel = 79;
			18192: Pixel = 107;
			18193: Pixel = 88;
			18194: Pixel = 135;
			18195: Pixel = 138;
			18196: Pixel = 120;
			18197: Pixel = 128;
			18198: Pixel = 94;
			18199: Pixel = 134;
			18200: Pixel = 104;
			18201: Pixel = 102;
			18202: Pixel = 93;
			18203: Pixel = 37;
			18204: Pixel = 48;
			18205: Pixel = 73;
			18206: Pixel = 62;
			18207: Pixel = 56;
			18208: Pixel = 52;
			18209: Pixel = 49;
			18210: Pixel = 55;
			18211: Pixel = 67;
			18212: Pixel = 58;
			18213: Pixel = 50;
			18214: Pixel = 61;
			18215: Pixel = 68;
			18216: Pixel = 82;
			18217: Pixel = 113;
			18218: Pixel = 70;
			18219: Pixel = 45;
			18220: Pixel = 86;
			18221: Pixel = 122;
			18222: Pixel = 115;
			18223: Pixel = 115;
			18224: Pixel = 126;
			18225: Pixel = 134;
			18226: Pixel = 137;
			18227: Pixel = 138;
			18228: Pixel = 139;
			18229: Pixel = 140;
			18230: Pixel = 139;
			18231: Pixel = 140;
			18232: Pixel = 142;
			18233: Pixel = 148;
			18234: Pixel = 152;
			18235: Pixel = 159;
			18236: Pixel = 161;
			18237: Pixel = 164;
			18238: Pixel = 168;
			18239: Pixel = 174;
			18240: Pixel = 175;
			18241: Pixel = 178;
			18242: Pixel = 183;
			18243: Pixel = 184;
			18244: Pixel = 192;
			18245: Pixel = 196;
			18246: Pixel = 201;
			18247: Pixel = 204;
			18248: Pixel = 208;
			18249: Pixel = 211;
			18250: Pixel = 211;
			18251: Pixel = 225;
			18252: Pixel = 179;
			18253: Pixel = 56;
			18254: Pixel = 43;
			18255: Pixel = 54;
			18256: Pixel = 67;
			18257: Pixel = 68;
			18258: Pixel = 45;
			18259: Pixel = 121;
			18260: Pixel = 151;
			18261: Pixel = 139;
			18262: Pixel = 149;
			18263: Pixel = 147;
			18264: Pixel = 145;
			18265: Pixel = 142;
			18266: Pixel = 142;
			18267: Pixel = 142;
			18268: Pixel = 141;
			18269: Pixel = 140;
			18270: Pixel = 138;
			18271: Pixel = 135;
			18272: Pixel = 133;
			18273: Pixel = 130;
			18274: Pixel = 127;
			18275: Pixel = 124;
			18276: Pixel = 121;
			18277: Pixel = 128;
			18278: Pixel = 135;
			18279: Pixel = 118;
			18280: Pixel = 150;
			18281: Pixel = 206;
			18282: Pixel = 212;
			18283: Pixel = 212;
			18284: Pixel = 213;
			18285: Pixel = 212;
			18286: Pixel = 200;
			18287: Pixel = 169;
			18288: Pixel = 100;
			18289: Pixel = 58;
			18290: Pixel = 89;
			18291: Pixel = 92;
			18292: Pixel = 91;
			18293: Pixel = 91;
			18294: Pixel = 100;
			18295: Pixel = 114;
			18296: Pixel = 106;
			18297: Pixel = 92;
			18298: Pixel = 89;
			18299: Pixel = 100;
			18300: Pixel = 57;
			18301: Pixel = 104;
			18302: Pixel = 135;
			18303: Pixel = 157;
			18304: Pixel = 165;
			18305: Pixel = 153;
			18306: Pixel = 119;
			18307: Pixel = 55;
			18308: Pixel = 57;
			18309: Pixel = 113;
			18310: Pixel = 151;
			18311: Pixel = 169;
			18312: Pixel = 178;
			18313: Pixel = 176;
			18314: Pixel = 177;
			18315: Pixel = 179;
			18316: Pixel = 171;
			18317: Pixel = 149;
			18318: Pixel = 166;
			18319: Pixel = 124;
			18320: Pixel = 61;
			18321: Pixel = 40;
			18322: Pixel = 43;
			18323: Pixel = 43;
			18324: Pixel = 43;
			18325: Pixel = 65;
			18326: Pixel = 57;
			18327: Pixel = 55;
			18328: Pixel = 49;
			18329: Pixel = 37;
			18330: Pixel = 85;
			18331: Pixel = 85;
			18332: Pixel = 64;
			18333: Pixel = 45;
			18334: Pixel = 55;
			18335: Pixel = 85;
			18336: Pixel = 34;
			18337: Pixel = 82;
			18338: Pixel = 88;
			18339: Pixel = 58;
			18340: Pixel = 75;
			18341: Pixel = 70;
			18342: Pixel = 88;
			18343: Pixel = 102;
			18344: Pixel = 121;
			18345: Pixel = 120;
			18346: Pixel = 132;
			18347: Pixel = 148;
			18348: Pixel = 129;
			18349: Pixel = 64;
			18350: Pixel = 125;
			18351: Pixel = 116;
			18352: Pixel = 125;
			18353: Pixel = 26;
			18354: Pixel = 41;
			18355: Pixel = 67;
			18356: Pixel = 61;
			18357: Pixel = 55;
			18358: Pixel = 50;
			18359: Pixel = 46;
			18360: Pixel = 52;
			18361: Pixel = 64;
			18362: Pixel = 55;
			18363: Pixel = 46;
			18364: Pixel = 53;
			18365: Pixel = 64;
			18366: Pixel = 91;
			18367: Pixel = 123;
			18368: Pixel = 82;
			18369: Pixel = 43;
			18370: Pixel = 82;
			18371: Pixel = 110;
			18372: Pixel = 113;
			18373: Pixel = 131;
			18374: Pixel = 133;
			18375: Pixel = 130;
			18376: Pixel = 137;
			18377: Pixel = 138;
			18378: Pixel = 140;
			18379: Pixel = 138;
			18380: Pixel = 138;
			18381: Pixel = 141;
			18382: Pixel = 143;
			18383: Pixel = 146;
			18384: Pixel = 150;
			18385: Pixel = 154;
			18386: Pixel = 160;
			18387: Pixel = 161;
			18388: Pixel = 165;
			18389: Pixel = 172;
			18390: Pixel = 173;
			18391: Pixel = 177;
			18392: Pixel = 181;
			18393: Pixel = 184;
			18394: Pixel = 190;
			18395: Pixel = 194;
			18396: Pixel = 197;
			18397: Pixel = 202;
			18398: Pixel = 206;
			18399: Pixel = 209;
			18400: Pixel = 213;
			18401: Pixel = 214;
			18402: Pixel = 229;
			18403: Pixel = 145;
			18404: Pixel = 38;
			18405: Pixel = 51;
			18406: Pixel = 58;
			18407: Pixel = 58;
			18408: Pixel = 44;
			18409: Pixel = 133;
			18410: Pixel = 145;
			18411: Pixel = 141;
			18412: Pixel = 147;
			18413: Pixel = 146;
			18414: Pixel = 145;
			18415: Pixel = 143;
			18416: Pixel = 144;
			18417: Pixel = 142;
			18418: Pixel = 142;
			18419: Pixel = 141;
			18420: Pixel = 140;
			18421: Pixel = 136;
			18422: Pixel = 135;
			18423: Pixel = 133;
			18424: Pixel = 127;
			18425: Pixel = 127;
			18426: Pixel = 126;
			18427: Pixel = 135;
			18428: Pixel = 137;
			18429: Pixel = 125;
			18430: Pixel = 168;
			18431: Pixel = 213;
			18432: Pixel = 214;
			18433: Pixel = 212;
			18434: Pixel = 212;
			18435: Pixel = 210;
			18436: Pixel = 194;
			18437: Pixel = 135;
			18438: Pixel = 76;
			18439: Pixel = 79;
			18440: Pixel = 96;
			18441: Pixel = 91;
			18442: Pixel = 94;
			18443: Pixel = 100;
			18444: Pixel = 113;
			18445: Pixel = 109;
			18446: Pixel = 96;
			18447: Pixel = 92;
			18448: Pixel = 99;
			18449: Pixel = 103;
			18450: Pixel = 38;
			18451: Pixel = 72;
			18452: Pixel = 123;
			18453: Pixel = 161;
			18454: Pixel = 168;
			18455: Pixel = 158;
			18456: Pixel = 132;
			18457: Pixel = 63;
			18458: Pixel = 49;
			18459: Pixel = 112;
			18460: Pixel = 153;
			18461: Pixel = 169;
			18462: Pixel = 177;
			18463: Pixel = 176;
			18464: Pixel = 177;
			18465: Pixel = 178;
			18466: Pixel = 170;
			18467: Pixel = 151;
			18468: Pixel = 152;
			18469: Pixel = 136;
			18470: Pixel = 87;
			18471: Pixel = 38;
			18472: Pixel = 43;
			18473: Pixel = 43;
			18474: Pixel = 53;
			18475: Pixel = 74;
			18476: Pixel = 45;
			18477: Pixel = 51;
			18478: Pixel = 53;
			18479: Pixel = 42;
			18480: Pixel = 98;
			18481: Pixel = 81;
			18482: Pixel = 58;
			18483: Pixel = 53;
			18484: Pixel = 34;
			18485: Pixel = 82;
			18486: Pixel = 61;
			18487: Pixel = 64;
			18488: Pixel = 73;
			18489: Pixel = 86;
			18490: Pixel = 83;
			18491: Pixel = 97;
			18492: Pixel = 73;
			18493: Pixel = 91;
			18494: Pixel = 103;
			18495: Pixel = 114;
			18496: Pixel = 119;
			18497: Pixel = 156;
			18498: Pixel = 149;
			18499: Pixel = 43;
			18500: Pixel = 64;
			18501: Pixel = 137;
			18502: Pixel = 145;
			18503: Pixel = 30;
			18504: Pixel = 38;
			18505: Pixel = 62;
			18506: Pixel = 63;
			18507: Pixel = 57;
			18508: Pixel = 49;
			18509: Pixel = 45;
			18510: Pixel = 52;
			18511: Pixel = 70;
			18512: Pixel = 56;
			18513: Pixel = 53;
			18514: Pixel = 51;
			18515: Pixel = 61;
			18516: Pixel = 101;
			18517: Pixel = 123;
			18518: Pixel = 89;
			18519: Pixel = 40;
			18520: Pixel = 75;
			18521: Pixel = 110;
			18522: Pixel = 123;
			18523: Pixel = 132;
			18524: Pixel = 132;
			18525: Pixel = 132;
			18526: Pixel = 134;
			18527: Pixel = 137;
			18528: Pixel = 140;
			18529: Pixel = 140;
			18530: Pixel = 141;
			18531: Pixel = 140;
			18532: Pixel = 142;
			18533: Pixel = 147;
			18534: Pixel = 150;
			18535: Pixel = 153;
			18536: Pixel = 158;
			18537: Pixel = 161;
			18538: Pixel = 164;
			18539: Pixel = 168;
			18540: Pixel = 171;
			18541: Pixel = 175;
			18542: Pixel = 181;
			18543: Pixel = 184;
			18544: Pixel = 189;
			18545: Pixel = 193;
			18546: Pixel = 196;
			18547: Pixel = 201;
			18548: Pixel = 204;
			18549: Pixel = 207;
			18550: Pixel = 211;
			18551: Pixel = 215;
			18552: Pixel = 221;
			18553: Pixel = 220;
			18554: Pixel = 81;
			18555: Pixel = 39;
			18556: Pixel = 56;
			18557: Pixel = 50;
			18558: Pixel = 47;
			18559: Pixel = 139;
			18560: Pixel = 139;
			18561: Pixel = 144;
			18562: Pixel = 147;
			18563: Pixel = 146;
			18564: Pixel = 144;
			18565: Pixel = 143;
			18566: Pixel = 144;
			18567: Pixel = 140;
			18568: Pixel = 140;
			18569: Pixel = 140;
			18570: Pixel = 138;
			18571: Pixel = 138;
			18572: Pixel = 137;
			18573: Pixel = 133;
			18574: Pixel = 128;
			18575: Pixel = 127;
			18576: Pixel = 123;
			18577: Pixel = 130;
			18578: Pixel = 143;
			18579: Pixel = 149;
			18580: Pixel = 184;
			18581: Pixel = 214;
			18582: Pixel = 214;
			18583: Pixel = 213;
			18584: Pixel = 210;
			18585: Pixel = 208;
			18586: Pixel = 181;
			18587: Pixel = 100;
			18588: Pixel = 74;
			18589: Pixel = 91;
			18590: Pixel = 90;
			18591: Pixel = 97;
			18592: Pixel = 101;
			18593: Pixel = 110;
			18594: Pixel = 110;
			18595: Pixel = 93;
			18596: Pixel = 89;
			18597: Pixel = 99;
			18598: Pixel = 104;
			18599: Pixel = 103;
			18600: Pixel = 34;
			18601: Pixel = 46;
			18602: Pixel = 111;
			18603: Pixel = 162;
			18604: Pixel = 170;
			18605: Pixel = 165;
			18606: Pixel = 140;
			18607: Pixel = 62;
			18608: Pixel = 39;
			18609: Pixel = 108;
			18610: Pixel = 152;
			18611: Pixel = 168;
			18612: Pixel = 177;
			18613: Pixel = 175;
			18614: Pixel = 175;
			18615: Pixel = 179;
			18616: Pixel = 172;
			18617: Pixel = 159;
			18618: Pixel = 124;
			18619: Pixel = 131;
			18620: Pixel = 76;
			18621: Pixel = 38;
			18622: Pixel = 46;
			18623: Pixel = 45;
			18624: Pixel = 62;
			18625: Pixel = 53;
			18626: Pixel = 44;
			18627: Pixel = 49;
			18628: Pixel = 44;
			18629: Pixel = 42;
			18630: Pixel = 106;
			18631: Pixel = 79;
			18632: Pixel = 57;
			18633: Pixel = 63;
			18634: Pixel = 34;
			18635: Pixel = 43;
			18636: Pixel = 78;
			18637: Pixel = 88;
			18638: Pixel = 67;
			18639: Pixel = 71;
			18640: Pixel = 87;
			18641: Pixel = 106;
			18642: Pixel = 110;
			18643: Pixel = 80;
			18644: Pixel = 85;
			18645: Pixel = 120;
			18646: Pixel = 140;
			18647: Pixel = 151;
			18648: Pixel = 107;
			18649: Pixel = 52;
			18650: Pixel = 58;
			18651: Pixel = 161;
			18652: Pixel = 162;
			18653: Pixel = 34;
			18654: Pixel = 38;
			18655: Pixel = 64;
			18656: Pixel = 66;
			18657: Pixel = 63;
			18658: Pixel = 46;
			18659: Pixel = 47;
			18660: Pixel = 53;
			18661: Pixel = 65;
			18662: Pixel = 50;
			18663: Pixel = 51;
			18664: Pixel = 50;
			18665: Pixel = 68;
			18666: Pixel = 106;
			18667: Pixel = 112;
			18668: Pixel = 89;
			18669: Pixel = 43;
			18670: Pixel = 77;
			18671: Pixel = 114;
			18672: Pixel = 123;
			18673: Pixel = 130;
			18674: Pixel = 128;
			18675: Pixel = 135;
			18676: Pixel = 133;
			18677: Pixel = 136;
			18678: Pixel = 138;
			18679: Pixel = 140;
			18680: Pixel = 140;
			18681: Pixel = 141;
			18682: Pixel = 146;
			18683: Pixel = 148;
			18684: Pixel = 148;
			18685: Pixel = 151;
			18686: Pixel = 155;
			18687: Pixel = 159;
			18688: Pixel = 162;
			18689: Pixel = 166;
			18690: Pixel = 171;
			18691: Pixel = 174;
			18692: Pixel = 179;
			18693: Pixel = 181;
			18694: Pixel = 187;
			18695: Pixel = 191;
			18696: Pixel = 196;
			18697: Pixel = 201;
			18698: Pixel = 205;
			18699: Pixel = 208;
			18700: Pixel = 211;
			18701: Pixel = 215;
			18702: Pixel = 216;
			18703: Pixel = 229;
			18704: Pixel = 164;
			18705: Pixel = 36;
			18706: Pixel = 47;
			18707: Pixel = 39;
			18708: Pixel = 51;
			18709: Pixel = 148;
			18710: Pixel = 140;
			18711: Pixel = 147;
			18712: Pixel = 148;
			18713: Pixel = 145;
			18714: Pixel = 145;
			18715: Pixel = 143;
			18716: Pixel = 144;
			18717: Pixel = 140;
			18718: Pixel = 140;
			18719: Pixel = 138;
			18720: Pixel = 136;
			18721: Pixel = 137;
			18722: Pixel = 134;
			18723: Pixel = 132;
			18724: Pixel = 126;
			18725: Pixel = 123;
			18726: Pixel = 121;
			18727: Pixel = 143;
			18728: Pixel = 172;
			18729: Pixel = 188;
			18730: Pixel = 201;
			18731: Pixel = 213;
			18732: Pixel = 215;
			18733: Pixel = 213;
			18734: Pixel = 209;
			18735: Pixel = 203;
			18736: Pixel = 153;
			18737: Pixel = 87;
			18738: Pixel = 89;
			18739: Pixel = 94;
			18740: Pixel = 91;
			18741: Pixel = 102;
			18742: Pixel = 109;
			18743: Pixel = 112;
			18744: Pixel = 97;
			18745: Pixel = 86;
			18746: Pixel = 91;
			18747: Pixel = 103;
			18748: Pixel = 102;
			18749: Pixel = 100;
			18750: Pixel = 35;
			18751: Pixel = 46;
			18752: Pixel = 100;
			18753: Pixel = 159;
			18754: Pixel = 173;
			18755: Pixel = 168;
			18756: Pixel = 139;
			18757: Pixel = 53;
			18758: Pixel = 41;
			18759: Pixel = 109;
			18760: Pixel = 151;
			18761: Pixel = 169;
			18762: Pixel = 180;
			18763: Pixel = 177;
			18764: Pixel = 177;
			18765: Pixel = 180;
			18766: Pixel = 174;
			18767: Pixel = 160;
			18768: Pixel = 131;
			18769: Pixel = 126;
			18770: Pixel = 84;
			18771: Pixel = 42;
			18772: Pixel = 45;
			18773: Pixel = 52;
			18774: Pixel = 55;
			18775: Pixel = 49;
			18776: Pixel = 47;
			18777: Pixel = 50;
			18778: Pixel = 49;
			18779: Pixel = 47;
			18780: Pixel = 129;
			18781: Pixel = 69;
			18782: Pixel = 46;
			18783: Pixel = 69;
			18784: Pixel = 42;
			18785: Pixel = 51;
			18786: Pixel = 54;
			18787: Pixel = 68;
			18788: Pixel = 62;
			18789: Pixel = 64;
			18790: Pixel = 81;
			18791: Pixel = 101;
			18792: Pixel = 99;
			18793: Pixel = 84;
			18794: Pixel = 79;
			18795: Pixel = 113;
			18796: Pixel = 149;
			18797: Pixel = 147;
			18798: Pixel = 123;
			18799: Pixel = 41;
			18800: Pixel = 52;
			18801: Pixel = 169;
			18802: Pixel = 141;
			18803: Pixel = 23;
			18804: Pixel = 44;
			18805: Pixel = 68;
			18806: Pixel = 70;
			18807: Pixel = 69;
			18808: Pixel = 48;
			18809: Pixel = 49;
			18810: Pixel = 52;
			18811: Pixel = 63;
			18812: Pixel = 45;
			18813: Pixel = 50;
			18814: Pixel = 54;
			18815: Pixel = 83;
			18816: Pixel = 106;
			18817: Pixel = 103;
			18818: Pixel = 99;
			18819: Pixel = 49;
			18820: Pixel = 78;
			18821: Pixel = 112;
			18822: Pixel = 128;
			18823: Pixel = 129;
			18824: Pixel = 128;
			18825: Pixel = 135;
			18826: Pixel = 138;
			18827: Pixel = 139;
			18828: Pixel = 136;
			18829: Pixel = 138;
			18830: Pixel = 139;
			18831: Pixel = 141;
			18832: Pixel = 144;
			18833: Pixel = 146;
			18834: Pixel = 146;
			18835: Pixel = 151;
			18836: Pixel = 155;
			18837: Pixel = 156;
			18838: Pixel = 160;
			18839: Pixel = 165;
			18840: Pixel = 170;
			18841: Pixel = 174;
			18842: Pixel = 176;
			18843: Pixel = 183;
			18844: Pixel = 186;
			18845: Pixel = 189;
			18846: Pixel = 195;
			18847: Pixel = 201;
			18848: Pixel = 206;
			18849: Pixel = 208;
			18850: Pixel = 211;
			18851: Pixel = 213;
			18852: Pixel = 217;
			18853: Pixel = 221;
			18854: Pixel = 219;
			18855: Pixel = 76;
			18856: Pixel = 32;
			18857: Pixel = 33;
			18858: Pixel = 59;
			18859: Pixel = 152;
			18860: Pixel = 141;
			18861: Pixel = 147;
			18862: Pixel = 149;
			18863: Pixel = 148;
			18864: Pixel = 145;
			18865: Pixel = 145;
			18866: Pixel = 143;
			18867: Pixel = 142;
			18868: Pixel = 139;
			18869: Pixel = 137;
			18870: Pixel = 134;
			18871: Pixel = 135;
			18872: Pixel = 133;
			18873: Pixel = 128;
			18874: Pixel = 124;
			18875: Pixel = 121;
			18876: Pixel = 139;
			18877: Pixel = 178;
			18878: Pixel = 195;
			18879: Pixel = 200;
			18880: Pixel = 208;
			18881: Pixel = 216;
			18882: Pixel = 215;
			18883: Pixel = 213;
			18884: Pixel = 208;
			18885: Pixel = 187;
			18886: Pixel = 118;
			18887: Pixel = 87;
			18888: Pixel = 94;
			18889: Pixel = 93;
			18890: Pixel = 100;
			18891: Pixel = 106;
			18892: Pixel = 113;
			18893: Pixel = 105;
			18894: Pixel = 91;
			18895: Pixel = 90;
			18896: Pixel = 99;
			18897: Pixel = 103;
			18898: Pixel = 98;
			18899: Pixel = 104;
			18900: Pixel = 32;
			18901: Pixel = 40;
			18902: Pixel = 94;
			18903: Pixel = 152;
			18904: Pixel = 169;
			18905: Pixel = 168;
			18906: Pixel = 136;
			18907: Pixel = 56;
			18908: Pixel = 38;
			18909: Pixel = 105;
			18910: Pixel = 151;
			18911: Pixel = 170;
			18912: Pixel = 178;
			18913: Pixel = 177;
			18914: Pixel = 177;
			18915: Pixel = 181;
			18916: Pixel = 176;
			18917: Pixel = 156;
			18918: Pixel = 147;
			18919: Pixel = 141;
			18920: Pixel = 59;
			18921: Pixel = 45;
			18922: Pixel = 47;
			18923: Pixel = 60;
			18924: Pixel = 46;
			18925: Pixel = 47;
			18926: Pixel = 43;
			18927: Pixel = 51;
			18928: Pixel = 35;
			18929: Pixel = 70;
			18930: Pixel = 140;
			18931: Pixel = 64;
			18932: Pixel = 40;
			18933: Pixel = 61;
			18934: Pixel = 52;
			18935: Pixel = 60;
			18936: Pixel = 55;
			18937: Pixel = 46;
			18938: Pixel = 45;
			18939: Pixel = 62;
			18940: Pixel = 76;
			18941: Pixel = 97;
			18942: Pixel = 109;
			18943: Pixel = 86;
			18944: Pixel = 67;
			18945: Pixel = 117;
			18946: Pixel = 134;
			18947: Pixel = 134;
			18948: Pixel = 137;
			18949: Pixel = 84;
			18950: Pixel = 45;
			18951: Pixel = 155;
			18952: Pixel = 107;
			18953: Pixel = 45;
			18954: Pixel = 43;
			18955: Pixel = 76;
			18956: Pixel = 67;
			18957: Pixel = 62;
			18958: Pixel = 52;
			18959: Pixel = 49;
			18960: Pixel = 52;
			18961: Pixel = 61;
			18962: Pixel = 52;
			18963: Pixel = 48;
			18964: Pixel = 59;
			18965: Pixel = 88;
			18966: Pixel = 105;
			18967: Pixel = 121;
			18968: Pixel = 107;
			18969: Pixel = 48;
			18970: Pixel = 83;
			18971: Pixel = 113;
			18972: Pixel = 131;
			18973: Pixel = 130;
			18974: Pixel = 132;
			18975: Pixel = 136;
			18976: Pixel = 136;
			18977: Pixel = 138;
			18978: Pixel = 136;
			18979: Pixel = 135;
			18980: Pixel = 137;
			18981: Pixel = 139;
			18982: Pixel = 144;
			18983: Pixel = 145;
			18984: Pixel = 145;
			18985: Pixel = 150;
			18986: Pixel = 153;
			18987: Pixel = 155;
			18988: Pixel = 159;
			18989: Pixel = 165;
			18990: Pixel = 167;
			18991: Pixel = 171;
			18992: Pixel = 176;
			18993: Pixel = 179;
			18994: Pixel = 185;
			18995: Pixel = 189;
			18996: Pixel = 194;
			18997: Pixel = 199;
			18998: Pixel = 204;
			18999: Pixel = 208;
			19000: Pixel = 210;
			19001: Pixel = 212;
			19002: Pixel = 215;
			19003: Pixel = 216;
			19004: Pixel = 232;
			19005: Pixel = 143;
			19006: Pixel = 29;
			19007: Pixel = 30;
			19008: Pixel = 73;
			19009: Pixel = 150;
			19010: Pixel = 143;
			19011: Pixel = 148;
			19012: Pixel = 147;
			19013: Pixel = 147;
			19014: Pixel = 146;
			19015: Pixel = 145;
			19016: Pixel = 142;
			19017: Pixel = 140;
			19018: Pixel = 139;
			19019: Pixel = 134;
			19020: Pixel = 133;
			19021: Pixel = 132;
			19022: Pixel = 129;
			19023: Pixel = 127;
			19024: Pixel = 124;
			19025: Pixel = 123;
			19026: Pixel = 173;
			19027: Pixel = 208;
			19028: Pixel = 207;
			19029: Pixel = 202;
			19030: Pixel = 209;
			19031: Pixel = 217;
			19032: Pixel = 215;
			19033: Pixel = 213;
			19034: Pixel = 203;
			19035: Pixel = 158;
			19036: Pixel = 98;
			19037: Pixel = 91;
			19038: Pixel = 92;
			19039: Pixel = 95;
			19040: Pixel = 106;
			19041: Pixel = 113;
			19042: Pixel = 115;
			19043: Pixel = 97;
			19044: Pixel = 88;
			19045: Pixel = 94;
			19046: Pixel = 104;
			19047: Pixel = 101;
			19048: Pixel = 100;
			19049: Pixel = 104;
			19050: Pixel = 31;
			19051: Pixel = 31;
			19052: Pixel = 82;
			19053: Pixel = 149;
			19054: Pixel = 170;
			19055: Pixel = 170;
			19056: Pixel = 142;
			19057: Pixel = 59;
			19058: Pixel = 36;
			19059: Pixel = 103;
			19060: Pixel = 152;
			19061: Pixel = 171;
			19062: Pixel = 179;
			19063: Pixel = 177;
			19064: Pixel = 178;
			19065: Pixel = 181;
			19066: Pixel = 174;
			19067: Pixel = 156;
			19068: Pixel = 145;
			19069: Pixel = 112;
			19070: Pixel = 40;
			19071: Pixel = 53;
			19072: Pixel = 57;
			19073: Pixel = 48;
			19074: Pixel = 43;
			19075: Pixel = 44;
			19076: Pixel = 47;
			19077: Pixel = 38;
			19078: Pixel = 42;
			19079: Pixel = 117;
			19080: Pixel = 120;
			19081: Pixel = 59;
			19082: Pixel = 38;
			19083: Pixel = 48;
			19084: Pixel = 60;
			19085: Pixel = 57;
			19086: Pixel = 44;
			19087: Pixel = 48;
			19088: Pixel = 53;
			19089: Pixel = 50;
			19090: Pixel = 67;
			19091: Pixel = 69;
			19092: Pixel = 121;
			19093: Pixel = 76;
			19094: Pixel = 54;
			19095: Pixel = 118;
			19096: Pixel = 143;
			19097: Pixel = 154;
			19098: Pixel = 109;
			19099: Pixel = 113;
			19100: Pixel = 111;
			19101: Pixel = 153;
			19102: Pixel = 153;
			19103: Pixel = 86;
			19104: Pixel = 39;
			19105: Pixel = 71;
			19106: Pixel = 59;
			19107: Pixel = 61;
			19108: Pixel = 56;
			19109: Pixel = 56;
			19110: Pixel = 51;
			19111: Pixel = 50;
			19112: Pixel = 54;
			19113: Pixel = 55;
			19114: Pixel = 71;
			19115: Pixel = 108;
			19116: Pixel = 123;
			19117: Pixel = 126;
			19118: Pixel = 105;
			19119: Pixel = 53;
			19120: Pixel = 88;
			19121: Pixel = 115;
			19122: Pixel = 129;
			19123: Pixel = 133;
			19124: Pixel = 136;
			19125: Pixel = 136;
			19126: Pixel = 137;
			19127: Pixel = 136;
			19128: Pixel = 135;
			19129: Pixel = 137;
			19130: Pixel = 136;
			19131: Pixel = 139;
			19132: Pixel = 143;
			19133: Pixel = 144;
			19134: Pixel = 145;
			19135: Pixel = 148;
			19136: Pixel = 151;
			19137: Pixel = 155;
			19138: Pixel = 159;
			19139: Pixel = 162;
			19140: Pixel = 163;
			19141: Pixel = 170;
			19142: Pixel = 175;
			19143: Pixel = 178;
			19144: Pixel = 184;
			19145: Pixel = 188;
			19146: Pixel = 193;
			19147: Pixel = 198;
			19148: Pixel = 204;
			19149: Pixel = 208;
			19150: Pixel = 209;
			19151: Pixel = 212;
			19152: Pixel = 214;
			19153: Pixel = 214;
			19154: Pixel = 226;
			19155: Pixel = 197;
			19156: Pixel = 42;
			19157: Pixel = 21;
			19158: Pixel = 86;
			19159: Pixel = 147;
			19160: Pixel = 146;
			19161: Pixel = 150;
			19162: Pixel = 146;
			19163: Pixel = 144;
			19164: Pixel = 144;
			19165: Pixel = 144;
			19166: Pixel = 141;
			19167: Pixel = 139;
			19168: Pixel = 139;
			19169: Pixel = 136;
			19170: Pixel = 133;
			19171: Pixel = 131;
			19172: Pixel = 126;
			19173: Pixel = 127;
			19174: Pixel = 120;
			19175: Pixel = 132;
			19176: Pixel = 198;
			19177: Pixel = 218;
			19178: Pixel = 214;
			19179: Pixel = 207;
			19180: Pixel = 211;
			19181: Pixel = 217;
			19182: Pixel = 216;
			19183: Pixel = 211;
			19184: Pixel = 186;
			19185: Pixel = 127;
			19186: Pixel = 94;
			19187: Pixel = 92;
			19188: Pixel = 89;
			19189: Pixel = 97;
			19190: Pixel = 108;
			19191: Pixel = 115;
			19192: Pixel = 107;
			19193: Pixel = 92;
			19194: Pixel = 89;
			19195: Pixel = 101;
			19196: Pixel = 105;
			19197: Pixel = 102;
			19198: Pixel = 103;
			19199: Pixel = 96;
			19200: Pixel = 31;
			19201: Pixel = 33;
			19202: Pixel = 77;
			19203: Pixel = 146;
			19204: Pixel = 172;
			19205: Pixel = 171;
			19206: Pixel = 145;
			19207: Pixel = 68;
			19208: Pixel = 34;
			19209: Pixel = 100;
			19210: Pixel = 151;
			19211: Pixel = 171;
			19212: Pixel = 178;
			19213: Pixel = 177;
			19214: Pixel = 179;
			19215: Pixel = 180;
			19216: Pixel = 175;
			19217: Pixel = 159;
			19218: Pixel = 141;
			19219: Pixel = 98;
			19220: Pixel = 53;
			19221: Pixel = 62;
			19222: Pixel = 46;
			19223: Pixel = 43;
			19224: Pixel = 45;
			19225: Pixel = 45;
			19226: Pixel = 44;
			19227: Pixel = 44;
			19228: Pixel = 96;
			19229: Pixel = 80;
			19230: Pixel = 93;
			19231: Pixel = 56;
			19232: Pixel = 40;
			19233: Pixel = 52;
			19234: Pixel = 71;
			19235: Pixel = 47;
			19236: Pixel = 44;
			19237: Pixel = 41;
			19238: Pixel = 63;
			19239: Pixel = 45;
			19240: Pixel = 66;
			19241: Pixel = 58;
			19242: Pixel = 108;
			19243: Pixel = 106;
			19244: Pixel = 93;
			19245: Pixel = 122;
			19246: Pixel = 145;
			19247: Pixel = 126;
			19248: Pixel = 128;
			19249: Pixel = 132;
			19250: Pixel = 169;
			19251: Pixel = 117;
			19252: Pixel = 48;
			19253: Pixel = 50;
			19254: Pixel = 56;
			19255: Pixel = 58;
			19256: Pixel = 56;
			19257: Pixel = 59;
			19258: Pixel = 54;
			19259: Pixel = 55;
			19260: Pixel = 56;
			19261: Pixel = 51;
			19262: Pixel = 51;
			19263: Pixel = 64;
			19264: Pixel = 88;
			19265: Pixel = 123;
			19266: Pixel = 124;
			19267: Pixel = 125;
			19268: Pixel = 95;
			19269: Pixel = 55;
			19270: Pixel = 93;
			19271: Pixel = 116;
			19272: Pixel = 128;
			19273: Pixel = 131;
			19274: Pixel = 135;
			19275: Pixel = 137;
			19276: Pixel = 138;
			19277: Pixel = 138;
			19278: Pixel = 136;
			19279: Pixel = 137;
			19280: Pixel = 139;
			19281: Pixel = 138;
			19282: Pixel = 141;
			19283: Pixel = 143;
			19284: Pixel = 145;
			19285: Pixel = 147;
			19286: Pixel = 150;
			19287: Pixel = 155;
			19288: Pixel = 157;
			19289: Pixel = 160;
			19290: Pixel = 163;
			19291: Pixel = 168;
			19292: Pixel = 174;
			19293: Pixel = 178;
			19294: Pixel = 182;
			19295: Pixel = 188;
			19296: Pixel = 193;
			19297: Pixel = 197;
			19298: Pixel = 201;
			19299: Pixel = 206;
			19300: Pixel = 207;
			19301: Pixel = 210;
			19302: Pixel = 212;
			19303: Pixel = 214;
			19304: Pixel = 218;
			19305: Pixel = 223;
			19306: Pixel = 83;
			19307: Pixel = 16;
			19308: Pixel = 98;
			19309: Pixel = 145;
			19310: Pixel = 146;
			19311: Pixel = 149;
			19312: Pixel = 144;
			19313: Pixel = 145;
			19314: Pixel = 144;
			19315: Pixel = 142;
			19316: Pixel = 139;
			19317: Pixel = 139;
			19318: Pixel = 140;
			19319: Pixel = 137;
			19320: Pixel = 132;
			19321: Pixel = 132;
			19322: Pixel = 127;
			19323: Pixel = 124;
			19324: Pixel = 118;
			19325: Pixel = 144;
			19326: Pixel = 206;
			19327: Pixel = 218;
			19328: Pixel = 211;
			19329: Pixel = 208;
			19330: Pixel = 214;
			19331: Pixel = 217;
			19332: Pixel = 214;
			19333: Pixel = 204;
			19334: Pixel = 163;
			19335: Pixel = 113;
			19336: Pixel = 102;
			19337: Pixel = 97;
			19338: Pixel = 93;
			19339: Pixel = 99;
			19340: Pixel = 114;
			19341: Pixel = 112;
			19342: Pixel = 99;
			19343: Pixel = 91;
			19344: Pixel = 96;
			19345: Pixel = 105;
			19346: Pixel = 104;
			19347: Pixel = 98;
			19348: Pixel = 95;
			19349: Pixel = 85;
			19350: Pixel = 31;
			19351: Pixel = 31;
			19352: Pixel = 75;
			19353: Pixel = 145;
			19354: Pixel = 169;
			19355: Pixel = 170;
			19356: Pixel = 147;
			19357: Pixel = 79;
			19358: Pixel = 37;
			19359: Pixel = 97;
			19360: Pixel = 151;
			19361: Pixel = 171;
			19362: Pixel = 176;
			19363: Pixel = 174;
			19364: Pixel = 172;
			19365: Pixel = 173;
			19366: Pixel = 170;
			19367: Pixel = 156;
			19368: Pixel = 140;
			19369: Pixel = 113;
			19370: Pixel = 62;
			19371: Pixel = 50;
			19372: Pixel = 43;
			19373: Pixel = 45;
			19374: Pixel = 47;
			19375: Pixel = 47;
			19376: Pixel = 59;
			19377: Pixel = 76;
			19378: Pixel = 50;
			19379: Pixel = 54;
			19380: Pixel = 98;
			19381: Pixel = 69;
			19382: Pixel = 41;
			19383: Pixel = 55;
			19384: Pixel = 67;
			19385: Pixel = 47;
			19386: Pixel = 44;
			19387: Pixel = 46;
			19388: Pixel = 62;
			19389: Pixel = 45;
			19390: Pixel = 79;
			19391: Pixel = 58;
			19392: Pixel = 51;
			19393: Pixel = 88;
			19394: Pixel = 135;
			19395: Pixel = 129;
			19396: Pixel = 139;
			19397: Pixel = 103;
			19398: Pixel = 88;
			19399: Pixel = 124;
			19400: Pixel = 147;
			19401: Pixel = 142;
			19402: Pixel = 102;
			19403: Pixel = 98;
			19404: Pixel = 77;
			19405: Pixel = 63;
			19406: Pixel = 55;
			19407: Pixel = 63;
			19408: Pixel = 66;
			19409: Pixel = 52;
			19410: Pixel = 56;
			19411: Pixel = 48;
			19412: Pixel = 53;
			19413: Pixel = 72;
			19414: Pixel = 97;
			19415: Pixel = 124;
			19416: Pixel = 124;
			19417: Pixel = 128;
			19418: Pixel = 89;
			19419: Pixel = 55;
			19420: Pixel = 99;
			19421: Pixel = 119;
			19422: Pixel = 131;
			19423: Pixel = 132;
			19424: Pixel = 133;
			19425: Pixel = 139;
			19426: Pixel = 142;
			19427: Pixel = 139;
			19428: Pixel = 137;
			19429: Pixel = 135;
			19430: Pixel = 135;
			19431: Pixel = 137;
			19432: Pixel = 139;
			19433: Pixel = 141;
			19434: Pixel = 142;
			19435: Pixel = 146;
			19436: Pixel = 148;
			19437: Pixel = 153;
			19438: Pixel = 156;
			19439: Pixel = 159;
			19440: Pixel = 162;
			19441: Pixel = 166;
			19442: Pixel = 170;
			19443: Pixel = 174;
			19444: Pixel = 182;
			19445: Pixel = 189;
			19446: Pixel = 191;
			19447: Pixel = 196;
			19448: Pixel = 202;
			19449: Pixel = 205;
			19450: Pixel = 206;
			19451: Pixel = 210;
			19452: Pixel = 212;
			19453: Pixel = 214;
			19454: Pixel = 214;
			19455: Pixel = 230;
			19456: Pixel = 133;
			19457: Pixel = 15;
			19458: Pixel = 106;
			19459: Pixel = 145;
			19460: Pixel = 145;
			19461: Pixel = 151;
			19462: Pixel = 142;
			19463: Pixel = 143;
			19464: Pixel = 142;
			19465: Pixel = 140;
			19466: Pixel = 139;
			19467: Pixel = 139;
			19468: Pixel = 139;
			19469: Pixel = 137;
			19470: Pixel = 134;
			19471: Pixel = 131;
			19472: Pixel = 127;
			19473: Pixel = 125;
			19474: Pixel = 122;
			19475: Pixel = 154;
			19476: Pixel = 209;
			19477: Pixel = 214;
			19478: Pixel = 205;
			19479: Pixel = 206;
			19480: Pixel = 215;
			19481: Pixel = 217;
			19482: Pixel = 212;
			19483: Pixel = 188;
			19484: Pixel = 138;
			19485: Pixel = 116;
			19486: Pixel = 107;
			19487: Pixel = 98;
			19488: Pixel = 98;
			19489: Pixel = 101;
			19490: Pixel = 112;
			19491: Pixel = 109;
			19492: Pixel = 96;
			19493: Pixel = 90;
			19494: Pixel = 99;
			19495: Pixel = 105;
			19496: Pixel = 102;
			19497: Pixel = 95;
			19498: Pixel = 88;
			19499: Pixel = 81;
			19500: Pixel = 30;
			19501: Pixel = 30;
			19502: Pixel = 67;
			19503: Pixel = 139;
			19504: Pixel = 170;
			19505: Pixel = 171;
			19506: Pixel = 154;
			19507: Pixel = 82;
			19508: Pixel = 37;
			19509: Pixel = 95;
			19510: Pixel = 149;
			19511: Pixel = 170;
			19512: Pixel = 177;
			19513: Pixel = 175;
			19514: Pixel = 173;
			19515: Pixel = 176;
			19516: Pixel = 172;
			19517: Pixel = 155;
			19518: Pixel = 145;
			19519: Pixel = 119;
			19520: Pixel = 60;
			19521: Pixel = 45;
			19522: Pixel = 47;
			19523: Pixel = 46;
			19524: Pixel = 48;
			19525: Pixel = 48;
			19526: Pixel = 56;
			19527: Pixel = 54;
			19528: Pixel = 47;
			19529: Pixel = 57;
			19530: Pixel = 85;
			19531: Pixel = 65;
			19532: Pixel = 49;
			19533: Pixel = 57;
			19534: Pixel = 50;
			19535: Pixel = 54;
			19536: Pixel = 48;
			19537: Pixel = 46;
			19538: Pixel = 58;
			19539: Pixel = 58;
			19540: Pixel = 87;
			19541: Pixel = 52;
			19542: Pixel = 36;
			19543: Pixel = 64;
			19544: Pixel = 128;
			19545: Pixel = 125;
			19546: Pixel = 124;
			19547: Pixel = 121;
			19548: Pixel = 74;
			19549: Pixel = 36;
			19550: Pixel = 74;
			19551: Pixel = 62;
			19552: Pixel = 91;
			19553: Pixel = 87;
			19554: Pixel = 108;
			19555: Pixel = 108;
			19556: Pixel = 120;
			19557: Pixel = 94;
			19558: Pixel = 63;
			19559: Pixel = 52;
			19560: Pixel = 54;
			19561: Pixel = 48;
			19562: Pixel = 61;
			19563: Pixel = 82;
			19564: Pixel = 109;
			19565: Pixel = 125;
			19566: Pixel = 125;
			19567: Pixel = 130;
			19568: Pixel = 84;
			19569: Pixel = 64;
			19570: Pixel = 104;
			19571: Pixel = 124;
			19572: Pixel = 131;
			19573: Pixel = 134;
			19574: Pixel = 133;
			19575: Pixel = 138;
			19576: Pixel = 141;
			19577: Pixel = 138;
			19578: Pixel = 138;
			19579: Pixel = 135;
			19580: Pixel = 133;
			19581: Pixel = 136;
			19582: Pixel = 138;
			19583: Pixel = 141;
			19584: Pixel = 142;
			19585: Pixel = 145;
			19586: Pixel = 150;
			19587: Pixel = 152;
			19588: Pixel = 154;
			19589: Pixel = 158;
			19590: Pixel = 158;
			19591: Pixel = 165;
			19592: Pixel = 168;
			19593: Pixel = 172;
			19594: Pixel = 180;
			19595: Pixel = 184;
			19596: Pixel = 190;
			19597: Pixel = 195;
			19598: Pixel = 199;
			19599: Pixel = 204;
			19600: Pixel = 206;
			19601: Pixel = 208;
			19602: Pixel = 211;
			19603: Pixel = 214;
			19604: Pixel = 213;
			19605: Pixel = 225;
			19606: Pixel = 178;
			19607: Pixel = 32;
			19608: Pixel = 113;
			19609: Pixel = 144;
			19610: Pixel = 143;
			19611: Pixel = 150;
			19612: Pixel = 146;
			19613: Pixel = 142;
			19614: Pixel = 142;
			19615: Pixel = 140;
			19616: Pixel = 138;
			19617: Pixel = 139;
			19618: Pixel = 139;
			19619: Pixel = 138;
			19620: Pixel = 135;
			19621: Pixel = 131;
			19622: Pixel = 125;
			19623: Pixel = 125;
			19624: Pixel = 124;
			19625: Pixel = 163;
			19626: Pixel = 210;
			19627: Pixel = 213;
			19628: Pixel = 203;
			19629: Pixel = 206;
			19630: Pixel = 217;
			19631: Pixel = 216;
			19632: Pixel = 206;
			19633: Pixel = 164;
			19634: Pixel = 120;
			19635: Pixel = 117;
			19636: Pixel = 107;
			19637: Pixel = 99;
			19638: Pixel = 97;
			19639: Pixel = 105;
			19640: Pixel = 109;
			19641: Pixel = 100;
			19642: Pixel = 88;
			19643: Pixel = 90;
			19644: Pixel = 103;
			19645: Pixel = 103;
			19646: Pixel = 95;
			19647: Pixel = 93;
			19648: Pixel = 88;
			19649: Pixel = 91;
			19650: Pixel = 33;
			19651: Pixel = 32;
			19652: Pixel = 57;
			19653: Pixel = 131;
			19654: Pixel = 166;
			19655: Pixel = 173;
			19656: Pixel = 157;
			19657: Pixel = 84;
			19658: Pixel = 40;
			19659: Pixel = 97;
			19660: Pixel = 148;
			19661: Pixel = 170;
			19662: Pixel = 176;
			19663: Pixel = 178;
			19664: Pixel = 178;
			19665: Pixel = 179;
			19666: Pixel = 175;
			19667: Pixel = 157;
			19668: Pixel = 149;
			19669: Pixel = 103;
			19670: Pixel = 48;
			19671: Pixel = 51;
			19672: Pixel = 50;
			19673: Pixel = 44;
			19674: Pixel = 48;
			19675: Pixel = 45;
			19676: Pixel = 45;
			19677: Pixel = 59;
			19678: Pixel = 52;
			19679: Pixel = 52;
			19680: Pixel = 71;
			19681: Pixel = 57;
			19682: Pixel = 55;
			19683: Pixel = 48;
			19684: Pixel = 54;
			19685: Pixel = 62;
			19686: Pixel = 40;
			19687: Pixel = 44;
			19688: Pixel = 51;
			19689: Pixel = 58;
			19690: Pixel = 88;
			19691: Pixel = 48;
			19692: Pixel = 74;
			19693: Pixel = 78;
			19694: Pixel = 105;
			19695: Pixel = 115;
			19696: Pixel = 112;
			19697: Pixel = 116;
			19698: Pixel = 135;
			19699: Pixel = 57;
			19700: Pixel = 72;
			19701: Pixel = 48;
			19702: Pixel = 41;
			19703: Pixel = 41;
			19704: Pixel = 59;
			19705: Pixel = 60;
			19706: Pixel = 72;
			19707: Pixel = 83;
			19708: Pixel = 84;
			19709: Pixel = 52;
			19710: Pixel = 48;
			19711: Pixel = 50;
			19712: Pixel = 74;
			19713: Pixel = 91;
			19714: Pixel = 116;
			19715: Pixel = 125;
			19716: Pixel = 129;
			19717: Pixel = 128;
			19718: Pixel = 73;
			19719: Pixel = 75;
			19720: Pixel = 110;
			19721: Pixel = 131;
			19722: Pixel = 132;
			19723: Pixel = 135;
			19724: Pixel = 138;
			19725: Pixel = 139;
			19726: Pixel = 139;
			19727: Pixel = 140;
			19728: Pixel = 139;
			19729: Pixel = 135;
			19730: Pixel = 134;
			19731: Pixel = 136;
			19732: Pixel = 138;
			19733: Pixel = 139;
			19734: Pixel = 141;
			19735: Pixel = 143;
			19736: Pixel = 146;
			19737: Pixel = 149;
			19738: Pixel = 154;
			19739: Pixel = 157;
			19740: Pixel = 158;
			19741: Pixel = 164;
			19742: Pixel = 167;
			19743: Pixel = 171;
			19744: Pixel = 175;
			19745: Pixel = 183;
			19746: Pixel = 190;
			19747: Pixel = 193;
			19748: Pixel = 197;
			19749: Pixel = 202;
			19750: Pixel = 206;
			19751: Pixel = 207;
			19752: Pixel = 210;
			19753: Pixel = 212;
			19754: Pixel = 213;
			19755: Pixel = 217;
			19756: Pixel = 208;
			19757: Pixel = 62;
			19758: Pixel = 114;
			19759: Pixel = 145;
			19760: Pixel = 147;
			19761: Pixel = 148;
			19762: Pixel = 144;
			19763: Pixel = 142;
			19764: Pixel = 144;
			19765: Pixel = 140;
			19766: Pixel = 139;
			19767: Pixel = 139;
			19768: Pixel = 140;
			19769: Pixel = 138;
			19770: Pixel = 135;
			19771: Pixel = 130;
			19772: Pixel = 128;
			19773: Pixel = 130;
			19774: Pixel = 126;
			19775: Pixel = 158;
			19776: Pixel = 204;
			19777: Pixel = 211;
			19778: Pixel = 202;
			19779: Pixel = 206;
			19780: Pixel = 219;
			19781: Pixel = 214;
			19782: Pixel = 196;
			19783: Pixel = 145;
			19784: Pixel = 116;
			19785: Pixel = 114;
			19786: Pixel = 108;
			19787: Pixel = 98;
			19788: Pixel = 93;
			19789: Pixel = 103;
			19790: Pixel = 100;
			19791: Pixel = 87;
			19792: Pixel = 87;
			19793: Pixel = 99;
			19794: Pixel = 105;
			19795: Pixel = 100;
			19796: Pixel = 95;
			19797: Pixel = 93;
			19798: Pixel = 90;
			19799: Pixel = 95;
			19800: Pixel = 37;
			19801: Pixel = 34;
			19802: Pixel = 52;
			19803: Pixel = 123;
			19804: Pixel = 163;
			19805: Pixel = 170;
			19806: Pixel = 155;
			19807: Pixel = 91;
			19808: Pixel = 46;
			19809: Pixel = 95;
			19810: Pixel = 146;
			19811: Pixel = 167;
			19812: Pixel = 176;
			19813: Pixel = 177;
			19814: Pixel = 177;
			19815: Pixel = 178;
			19816: Pixel = 175;
			19817: Pixel = 155;
			19818: Pixel = 153;
			19819: Pixel = 118;
			19820: Pixel = 55;
			19821: Pixel = 51;
			19822: Pixel = 46;
			19823: Pixel = 38;
			19824: Pixel = 46;
			19825: Pixel = 53;
			19826: Pixel = 74;
			19827: Pixel = 63;
			19828: Pixel = 45;
			19829: Pixel = 52;
			19830: Pixel = 62;
			19831: Pixel = 60;
			19832: Pixel = 54;
			19833: Pixel = 47;
			19834: Pixel = 50;
			19835: Pixel = 66;
			19836: Pixel = 41;
			19837: Pixel = 51;
			19838: Pixel = 49;
			19839: Pixel = 70;
			19840: Pixel = 75;
			19841: Pixel = 80;
			19842: Pixel = 65;
			19843: Pixel = 104;
			19844: Pixel = 97;
			19845: Pixel = 120;
			19846: Pixel = 114;
			19847: Pixel = 81;
			19848: Pixel = 121;
			19849: Pixel = 117;
			19850: Pixel = 75;
			19851: Pixel = 58;
			19852: Pixel = 41;
			19853: Pixel = 61;
			19854: Pixel = 54;
			19855: Pixel = 53;
			19856: Pixel = 59;
			19857: Pixel = 48;
			19858: Pixel = 59;
			19859: Pixel = 52;
			19860: Pixel = 43;
			19861: Pixel = 57;
			19862: Pixel = 81;
			19863: Pixel = 100;
			19864: Pixel = 117;
			19865: Pixel = 125;
			19866: Pixel = 129;
			19867: Pixel = 118;
			19868: Pixel = 62;
			19869: Pixel = 85;
			19870: Pixel = 117;
			19871: Pixel = 131;
			19872: Pixel = 134;
			19873: Pixel = 139;
			19874: Pixel = 138;
			19875: Pixel = 139;
			19876: Pixel = 141;
			19877: Pixel = 141;
			19878: Pixel = 140;
			19879: Pixel = 136;
			19880: Pixel = 136;
			19881: Pixel = 136;
			19882: Pixel = 138;
			19883: Pixel = 138;
			19884: Pixel = 140;
			19885: Pixel = 143;
			19886: Pixel = 147;
			19887: Pixel = 148;
			19888: Pixel = 153;
			19889: Pixel = 155;
			19890: Pixel = 159;
			19891: Pixel = 163;
			19892: Pixel = 166;
			19893: Pixel = 167;
			19894: Pixel = 174;
			19895: Pixel = 181;
			19896: Pixel = 187;
			19897: Pixel = 193;
			19898: Pixel = 197;
			19899: Pixel = 200;
			19900: Pixel = 204;
			19901: Pixel = 206;
			19902: Pixel = 208;
			19903: Pixel = 211;
			19904: Pixel = 212;
			19905: Pixel = 212;
			19906: Pixel = 221;
			19907: Pixel = 112;
			19908: Pixel = 112;
			19909: Pixel = 147;
			19910: Pixel = 145;
			19911: Pixel = 148;
			19912: Pixel = 144;
			19913: Pixel = 143;
			19914: Pixel = 143;
			19915: Pixel = 143;
			19916: Pixel = 142;
			19917: Pixel = 141;
			19918: Pixel = 141;
			19919: Pixel = 139;
			19920: Pixel = 136;
			19921: Pixel = 130;
			19922: Pixel = 130;
			19923: Pixel = 133;
			19924: Pixel = 133;
			19925: Pixel = 140;
			19926: Pixel = 175;
			19927: Pixel = 193;
			19928: Pixel = 193;
			19929: Pixel = 208;
			19930: Pixel = 218;
			19931: Pixel = 211;
			19932: Pixel = 187;
			19933: Pixel = 133;
			19934: Pixel = 112;
			19935: Pixel = 111;
			19936: Pixel = 104;
			19937: Pixel = 94;
			19938: Pixel = 94;
			19939: Pixel = 102;
			19940: Pixel = 83;
			19941: Pixel = 76;
			19942: Pixel = 101;
			19943: Pixel = 105;
			19944: Pixel = 100;
			19945: Pixel = 92;
			19946: Pixel = 93;
			19947: Pixel = 94;
			19948: Pixel = 94;
			19949: Pixel = 95;
			19950: Pixel = 41;
			19951: Pixel = 35;
			19952: Pixel = 44;
			19953: Pixel = 112;
			19954: Pixel = 162;
			19955: Pixel = 171;
			19956: Pixel = 157;
			19957: Pixel = 105;
			19958: Pixel = 54;
			19959: Pixel = 93;
			19960: Pixel = 146;
			19961: Pixel = 168;
			19962: Pixel = 176;
			19963: Pixel = 175;
			19964: Pixel = 176;
			19965: Pixel = 178;
			19966: Pixel = 173;
			19967: Pixel = 153;
			19968: Pixel = 155;
			19969: Pixel = 126;
			19970: Pixel = 71;
			19971: Pixel = 57;
			19972: Pixel = 38;
			19973: Pixel = 44;
			19974: Pixel = 67;
			19975: Pixel = 77;
			19976: Pixel = 61;
			19977: Pixel = 44;
			19978: Pixel = 43;
			19979: Pixel = 59;
			19980: Pixel = 65;
			19981: Pixel = 51;
			19982: Pixel = 53;
			19983: Pixel = 65;
			19984: Pixel = 52;
			19985: Pixel = 56;
			19986: Pixel = 61;
			19987: Pixel = 46;
			19988: Pixel = 68;
			19989: Pixel = 71;
			19990: Pixel = 50;
			19991: Pixel = 87;
			19992: Pixel = 56;
			19993: Pixel = 77;
			19994: Pixel = 122;
			19995: Pixel = 123;
			19996: Pixel = 118;
			19997: Pixel = 65;
			19998: Pixel = 69;
			19999: Pixel = 134;
			20000: Pixel = 127;
			20001: Pixel = 125;
			20002: Pixel = 54;
			20003: Pixel = 52;
			20004: Pixel = 50;
			20005: Pixel = 55;
			20006: Pixel = 56;
			20007: Pixel = 50;
			20008: Pixel = 49;
			20009: Pixel = 47;
			20010: Pixel = 45;
			20011: Pixel = 68;
			20012: Pixel = 89;
			20013: Pixel = 108;
			20014: Pixel = 120;
			20015: Pixel = 124;
			20016: Pixel = 127;
			20017: Pixel = 100;
			20018: Pixel = 59;
			20019: Pixel = 96;
			20020: Pixel = 122;
			20021: Pixel = 134;
			20022: Pixel = 137;
			20023: Pixel = 141;
			20024: Pixel = 140;
			20025: Pixel = 143;
			20026: Pixel = 142;
			20027: Pixel = 137;
			20028: Pixel = 138;
			20029: Pixel = 137;
			20030: Pixel = 136;
			20031: Pixel = 136;
			20032: Pixel = 135;
			20033: Pixel = 136;
			20034: Pixel = 141;
			20035: Pixel = 143;
			20036: Pixel = 146;
			20037: Pixel = 148;
			20038: Pixel = 151;
			20039: Pixel = 153;
			20040: Pixel = 156;
			20041: Pixel = 159;
			20042: Pixel = 163;
			20043: Pixel = 167;
			20044: Pixel = 172;
			20045: Pixel = 178;
			20046: Pixel = 184;
			20047: Pixel = 190;
			20048: Pixel = 195;
			20049: Pixel = 199;
			20050: Pixel = 202;
			20051: Pixel = 207;
			20052: Pixel = 209;
			20053: Pixel = 211;
			20054: Pixel = 212;
			20055: Pixel = 211;
			20056: Pixel = 221;
			20057: Pixel = 167;
			20058: Pixel = 125;
			20059: Pixel = 141;
			20060: Pixel = 122;
			20061: Pixel = 133;
			20062: Pixel = 136;
			20063: Pixel = 140;
			20064: Pixel = 144;
			20065: Pixel = 146;
			20066: Pixel = 145;
			20067: Pixel = 142;
			20068: Pixel = 143;
			20069: Pixel = 140;
			20070: Pixel = 137;
			20071: Pixel = 135;
			20072: Pixel = 135;
			20073: Pixel = 138;
			20074: Pixel = 141;
			20075: Pixel = 138;
			20076: Pixel = 138;
			20077: Pixel = 149;
			20078: Pixel = 179;
			20079: Pixel = 213;
			20080: Pixel = 217;
			20081: Pixel = 209;
			20082: Pixel = 177;
			20083: Pixel = 124;
			20084: Pixel = 109;
			20085: Pixel = 104;
			20086: Pixel = 94;
			20087: Pixel = 91;
			20088: Pixel = 100;
			20089: Pixel = 92;
			20090: Pixel = 76;
			20091: Pixel = 88;
			20092: Pixel = 108;
			20093: Pixel = 102;
			20094: Pixel = 93;
			20095: Pixel = 87;
			20096: Pixel = 92;
			20097: Pixel = 95;
			20098: Pixel = 97;
			20099: Pixel = 86;
			20100: Pixel = 38;
			20101: Pixel = 35;
			20102: Pixel = 42;
			20103: Pixel = 108;
			20104: Pixel = 158;
			20105: Pixel = 164;
			20106: Pixel = 155;
			20107: Pixel = 110;
			20108: Pixel = 58;
			20109: Pixel = 91;
			20110: Pixel = 143;
			20111: Pixel = 165;
			20112: Pixel = 175;
			20113: Pixel = 175;
			20114: Pixel = 175;
			20115: Pixel = 177;
			20116: Pixel = 174;
			20117: Pixel = 157;
			20118: Pixel = 145;
			20119: Pixel = 128;
			20120: Pixel = 74;
			20121: Pixel = 59;
			20122: Pixel = 42;
			20123: Pixel = 49;
			20124: Pixel = 59;
			20125: Pixel = 51;
			20126: Pixel = 44;
			20127: Pixel = 48;
			20128: Pixel = 48;
			20129: Pixel = 60;
			20130: Pixel = 65;
			20131: Pixel = 55;
			20132: Pixel = 66;
			20133: Pixel = 58;
			20134: Pixel = 56;
			20135: Pixel = 57;
			20136: Pixel = 56;
			20137: Pixel = 37;
			20138: Pixel = 81;
			20139: Pixel = 59;
			20140: Pixel = 36;
			20141: Pixel = 92;
			20142: Pixel = 96;
			20143: Pixel = 50;
			20144: Pixel = 49;
			20145: Pixel = 61;
			20146: Pixel = 124;
			20147: Pixel = 78;
			20148: Pixel = 55;
			20149: Pixel = 91;
			20150: Pixel = 155;
			20151: Pixel = 118;
			20152: Pixel = 39;
			20153: Pixel = 54;
			20154: Pixel = 44;
			20155: Pixel = 57;
			20156: Pixel = 49;
			20157: Pixel = 48;
			20158: Pixel = 44;
			20159: Pixel = 46;
			20160: Pixel = 51;
			20161: Pixel = 73;
			20162: Pixel = 99;
			20163: Pixel = 115;
			20164: Pixel = 120;
			20165: Pixel = 125;
			20166: Pixel = 125;
			20167: Pixel = 75;
			20168: Pixel = 66;
			20169: Pixel = 109;
			20170: Pixel = 131;
			20171: Pixel = 135;
			20172: Pixel = 137;
			20173: Pixel = 139;
			20174: Pixel = 140;
			20175: Pixel = 142;
			20176: Pixel = 145;
			20177: Pixel = 140;
			20178: Pixel = 140;
			20179: Pixel = 141;
			20180: Pixel = 138;
			20181: Pixel = 135;
			20182: Pixel = 138;
			20183: Pixel = 139;
			20184: Pixel = 141;
			20185: Pixel = 142;
			20186: Pixel = 146;
			20187: Pixel = 148;
			20188: Pixel = 149;
			20189: Pixel = 151;
			20190: Pixel = 154;
			20191: Pixel = 157;
			20192: Pixel = 160;
			20193: Pixel = 165;
			20194: Pixel = 172;
			20195: Pixel = 176;
			20196: Pixel = 181;
			20197: Pixel = 188;
			20198: Pixel = 194;
			20199: Pixel = 198;
			20200: Pixel = 201;
			20201: Pixel = 206;
			20202: Pixel = 210;
			20203: Pixel = 211;
			20204: Pixel = 212;
			20205: Pixel = 212;
			20206: Pixel = 216;
			20207: Pixel = 200;
			20208: Pixel = 141;
			20209: Pixel = 118;
			20210: Pixel = 94;
			20211: Pixel = 106;
			20212: Pixel = 111;
			20213: Pixel = 120;
			20214: Pixel = 130;
			20215: Pixel = 137;
			20216: Pixel = 142;
			20217: Pixel = 145;
			20218: Pixel = 144;
			20219: Pixel = 142;
			20220: Pixel = 140;
			20221: Pixel = 138;
			20222: Pixel = 140;
			20223: Pixel = 147;
			20224: Pixel = 147;
			20225: Pixel = 144;
			20226: Pixel = 135;
			20227: Pixel = 137;
			20228: Pixel = 183;
			20229: Pixel = 218;
			20230: Pixel = 218;
			20231: Pixel = 204;
			20232: Pixel = 159;
			20233: Pixel = 116;
			20234: Pixel = 109;
			20235: Pixel = 99;
			20236: Pixel = 89;
			20237: Pixel = 97;
			20238: Pixel = 95;
			20239: Pixel = 78;
			20240: Pixel = 81;
			20241: Pixel = 100;
			20242: Pixel = 103;
			20243: Pixel = 97;
			20244: Pixel = 89;
			20245: Pixel = 90;
			20246: Pixel = 96;
			20247: Pixel = 95;
			20248: Pixel = 91;
			20249: Pixel = 70;
			20250: Pixel = 36;
			20251: Pixel = 34;
			20252: Pixel = 42;
			20253: Pixel = 104;
			20254: Pixel = 156;
			20255: Pixel = 171;
			20256: Pixel = 163;
			20257: Pixel = 111;
			20258: Pixel = 59;
			20259: Pixel = 89;
			20260: Pixel = 141;
			20261: Pixel = 164;
			20262: Pixel = 173;
			20263: Pixel = 175;
			20264: Pixel = 176;
			20265: Pixel = 179;
			20266: Pixel = 174;
			20267: Pixel = 160;
			20268: Pixel = 138;
			20269: Pixel = 115;
			20270: Pixel = 79;
			20271: Pixel = 61;
			20272: Pixel = 40;
			20273: Pixel = 49;
			20274: Pixel = 50;
			20275: Pixel = 49;
			20276: Pixel = 46;
			20277: Pixel = 48;
			20278: Pixel = 59;
			20279: Pixel = 61;
			20280: Pixel = 57;
			20281: Pixel = 54;
			20282: Pixel = 77;
			20283: Pixel = 53;
			20284: Pixel = 42;
			20285: Pixel = 51;
			20286: Pixel = 43;
			20287: Pixel = 44;
			20288: Pixel = 64;
			20289: Pixel = 51;
			20290: Pixel = 60;
			20291: Pixel = 92;
			20292: Pixel = 129;
			20293: Pixel = 74;
			20294: Pixel = 54;
			20295: Pixel = 39;
			20296: Pixel = 76;
			20297: Pixel = 70;
			20298: Pixel = 66;
			20299: Pixel = 101;
			20300: Pixel = 108;
			20301: Pixel = 66;
			20302: Pixel = 44;
			20303: Pixel = 51;
			20304: Pixel = 44;
			20305: Pixel = 50;
			20306: Pixel = 47;
			20307: Pixel = 41;
			20308: Pixel = 40;
			20309: Pixel = 53;
			20310: Pixel = 64;
			20311: Pixel = 82;
			20312: Pixel = 108;
			20313: Pixel = 115;
			20314: Pixel = 120;
			20315: Pixel = 127;
			20316: Pixel = 111;
			20317: Pixel = 56;
			20318: Pixel = 79;
			20319: Pixel = 122;
			20320: Pixel = 135;
			20321: Pixel = 134;
			20322: Pixel = 137;
			20323: Pixel = 140;
			20324: Pixel = 141;
			20325: Pixel = 143;
			20326: Pixel = 143;
			20327: Pixel = 142;
			20328: Pixel = 141;
			20329: Pixel = 142;
			20330: Pixel = 139;
			20331: Pixel = 136;
			20332: Pixel = 136;
			20333: Pixel = 137;
			20334: Pixel = 139;
			20335: Pixel = 142;
			20336: Pixel = 146;
			20337: Pixel = 148;
			20338: Pixel = 149;
			20339: Pixel = 153;
			20340: Pixel = 152;
			20341: Pixel = 158;
			20342: Pixel = 161;
			20343: Pixel = 164;
			20344: Pixel = 168;
			20345: Pixel = 171;
			20346: Pixel = 178;
			20347: Pixel = 187;
			20348: Pixel = 191;
			20349: Pixel = 195;
			20350: Pixel = 201;
			20351: Pixel = 205;
			20352: Pixel = 209;
			20353: Pixel = 211;
			20354: Pixel = 213;
			20355: Pixel = 213;
			20356: Pixel = 214;
			20357: Pixel = 220;
			20358: Pixel = 144;
			20359: Pixel = 79;
			20360: Pixel = 75;
			20361: Pixel = 80;
			20362: Pixel = 83;
			20363: Pixel = 94;
			20364: Pixel = 102;
			20365: Pixel = 110;
			20366: Pixel = 120;
			20367: Pixel = 125;
			20368: Pixel = 132;
			20369: Pixel = 134;
			20370: Pixel = 138;
			20371: Pixel = 141;
			20372: Pixel = 147;
			20373: Pixel = 155;
			20374: Pixel = 148;
			20375: Pixel = 133;
			20376: Pixel = 130;
			20377: Pixel = 150;
			20378: Pixel = 198;
			20379: Pixel = 219;
			20380: Pixel = 215;
			20381: Pixel = 192;
			20382: Pixel = 141;
			20383: Pixel = 110;
			20384: Pixel = 95;
			20385: Pixel = 80;
			20386: Pixel = 88;
			20387: Pixel = 99;
			20388: Pixel = 80;
			20389: Pixel = 71;
			20390: Pixel = 94;
			20391: Pixel = 103;
			20392: Pixel = 96;
			20393: Pixel = 95;
			20394: Pixel = 89;
			20395: Pixel = 99;
			20396: Pixel = 101;
			20397: Pixel = 91;
			20398: Pixel = 79;
			20399: Pixel = 59;
			20400: Pixel = 34;
			20401: Pixel = 34;
			20402: Pixel = 38;
			20403: Pixel = 89;
			20404: Pixel = 164;
			20405: Pixel = 176;
			20406: Pixel = 169;
			20407: Pixel = 126;
			20408: Pixel = 60;
			20409: Pixel = 84;
			20410: Pixel = 139;
			20411: Pixel = 162;
			20412: Pixel = 172;
			20413: Pixel = 174;
			20414: Pixel = 176;
			20415: Pixel = 178;
			20416: Pixel = 175;
			20417: Pixel = 162;
			20418: Pixel = 141;
			20419: Pixel = 109;
			20420: Pixel = 86;
			20421: Pixel = 67;
			20422: Pixel = 37;
			20423: Pixel = 57;
			20424: Pixel = 47;
			20425: Pixel = 45;
			20426: Pixel = 44;
			20427: Pixel = 59;
			20428: Pixel = 58;
			20429: Pixel = 58;
			20430: Pixel = 54;
			20431: Pixel = 55;
			20432: Pixel = 68;
			20433: Pixel = 58;
			20434: Pixel = 47;
			20435: Pixel = 43;
			20436: Pixel = 48;
			20437: Pixel = 47;
			20438: Pixel = 51;
			20439: Pixel = 64;
			20440: Pixel = 81;
			20441: Pixel = 102;
			20442: Pixel = 123;
			20443: Pixel = 122;
			20444: Pixel = 63;
			20445: Pixel = 61;
			20446: Pixel = 61;
			20447: Pixel = 59;
			20448: Pixel = 94;
			20449: Pixel = 86;
			20450: Pixel = 85;
			20451: Pixel = 53;
			20452: Pixel = 47;
			20453: Pixel = 42;
			20454: Pixel = 49;
			20455: Pixel = 45;
			20456: Pixel = 46;
			20457: Pixel = 40;
			20458: Pixel = 45;
			20459: Pixel = 59;
			20460: Pixel = 76;
			20461: Pixel = 97;
			20462: Pixel = 118;
			20463: Pixel = 117;
			20464: Pixel = 117;
			20465: Pixel = 124;
			20466: Pixel = 73;
			20467: Pixel = 54;
			20468: Pixel = 101;
			20469: Pixel = 129;
			20470: Pixel = 133;
			20471: Pixel = 134;
			20472: Pixel = 135;
			20473: Pixel = 141;
			20474: Pixel = 142;
			20475: Pixel = 144;
			20476: Pixel = 141;
			20477: Pixel = 139;
			20478: Pixel = 142;
			20479: Pixel = 140;
			20480: Pixel = 139;
			20481: Pixel = 136;
			20482: Pixel = 136;
			20483: Pixel = 135;
			20484: Pixel = 137;
			20485: Pixel = 140;
			20486: Pixel = 143;
			20487: Pixel = 144;
			20488: Pixel = 148;
			20489: Pixel = 149;
			20490: Pixel = 153;
			20491: Pixel = 156;
			20492: Pixel = 159;
			20493: Pixel = 163;
			20494: Pixel = 169;
			20495: Pixel = 171;
			20496: Pixel = 174;
			20497: Pixel = 185;
			20498: Pixel = 188;
			20499: Pixel = 193;
			20500: Pixel = 200;
			20501: Pixel = 205;
			20502: Pixel = 207;
			20503: Pixel = 210;
			20504: Pixel = 212;
			20505: Pixel = 213;
			20506: Pixel = 214;
			20507: Pixel = 227;
			20508: Pixel = 154;
			20509: Pixel = 69;
			20510: Pixel = 84;
			20511: Pixel = 77;
			20512: Pixel = 73;
			20513: Pixel = 77;
			20514: Pixel = 78;
			20515: Pixel = 83;
			20516: Pixel = 87;
			20517: Pixel = 91;
			20518: Pixel = 99;
			20519: Pixel = 106;
			20520: Pixel = 115;
			20521: Pixel = 131;
			20522: Pixel = 149;
			20523: Pixel = 161;
			20524: Pixel = 147;
			20525: Pixel = 138;
			20526: Pixel = 135;
			20527: Pixel = 162;
			20528: Pixel = 211;
			20529: Pixel = 220;
			20530: Pixel = 208;
			20531: Pixel = 168;
			20532: Pixel = 122;
			20533: Pixel = 94;
			20534: Pixel = 77;
			20535: Pixel = 77;
			20536: Pixel = 95;
			20537: Pixel = 90;
			20538: Pixel = 71;
			20539: Pixel = 88;
			20540: Pixel = 104;
			20541: Pixel = 96;
			20542: Pixel = 93;
			20543: Pixel = 92;
			20544: Pixel = 94;
			20545: Pixel = 102;
			20546: Pixel = 99;
			20547: Pixel = 88;
			20548: Pixel = 67;
			20549: Pixel = 53;
			20550: Pixel = 38;
			20551: Pixel = 32;
			20552: Pixel = 30;
			20553: Pixel = 88;
			20554: Pixel = 162;
			20555: Pixel = 175;
			20556: Pixel = 171;
			20557: Pixel = 138;
			20558: Pixel = 68;
			20559: Pixel = 82;
			20560: Pixel = 137;
			20561: Pixel = 162;
			20562: Pixel = 171;
			20563: Pixel = 175;
			20564: Pixel = 176;
			20565: Pixel = 178;
			20566: Pixel = 176;
			20567: Pixel = 165;
			20568: Pixel = 126;
			20569: Pixel = 103;
			20570: Pixel = 95;
			20571: Pixel = 63;
			20572: Pixel = 42;
			20573: Pixel = 49;
			20574: Pixel = 42;
			20575: Pixel = 41;
			20576: Pixel = 56;
			20577: Pixel = 65;
			20578: Pixel = 46;
			20579: Pixel = 63;
			20580: Pixel = 50;
			20581: Pixel = 54;
			20582: Pixel = 66;
			20583: Pixel = 62;
			20584: Pixel = 59;
			20585: Pixel = 43;
			20586: Pixel = 49;
			20587: Pixel = 54;
			20588: Pixel = 53;
			20589: Pixel = 48;
			20590: Pixel = 43;
			20591: Pixel = 83;
			20592: Pixel = 106;
			20593: Pixel = 136;
			20594: Pixel = 126;
			20595: Pixel = 77;
			20596: Pixel = 97;
			20597: Pixel = 109;
			20598: Pixel = 77;
			20599: Pixel = 45;
			20600: Pixel = 43;
			20601: Pixel = 56;
			20602: Pixel = 50;
			20603: Pixel = 43;
			20604: Pixel = 46;
			20605: Pixel = 41;
			20606: Pixel = 43;
			20607: Pixel = 42;
			20608: Pixel = 48;
			20609: Pixel = 66;
			20610: Pixel = 86;
			20611: Pixel = 109;
			20612: Pixel = 119;
			20613: Pixel = 117;
			20614: Pixel = 123;
			20615: Pixel = 97;
			20616: Pixel = 40;
			20617: Pixel = 76;
			20618: Pixel = 120;
			20619: Pixel = 134;
			20620: Pixel = 134;
			20621: Pixel = 134;
			20622: Pixel = 136;
			20623: Pixel = 139;
			20624: Pixel = 140;
			20625: Pixel = 141;
			20626: Pixel = 141;
			20627: Pixel = 141;
			20628: Pixel = 142;
			20629: Pixel = 139;
			20630: Pixel = 139;
			20631: Pixel = 138;
			20632: Pixel = 136;
			20633: Pixel = 134;
			20634: Pixel = 136;
			20635: Pixel = 140;
			20636: Pixel = 141;
			20637: Pixel = 144;
			20638: Pixel = 145;
			20639: Pixel = 148;
			20640: Pixel = 150;
			20641: Pixel = 153;
			20642: Pixel = 158;
			20643: Pixel = 161;
			20644: Pixel = 166;
			20645: Pixel = 168;
			20646: Pixel = 173;
			20647: Pixel = 181;
			20648: Pixel = 187;
			20649: Pixel = 192;
			20650: Pixel = 199;
			20651: Pixel = 202;
			20652: Pixel = 206;
			20653: Pixel = 208;
			20654: Pixel = 211;
			20655: Pixel = 212;
			20656: Pixel = 213;
			20657: Pixel = 224;
			20658: Pixel = 185;
			20659: Pixel = 76;
			20660: Pixel = 92;
			20661: Pixel = 94;
			20662: Pixel = 88;
			20663: Pixel = 85;
			20664: Pixel = 78;
			20665: Pixel = 72;
			20666: Pixel = 66;
			20667: Pixel = 65;
			20668: Pixel = 65;
			20669: Pixel = 65;
			20670: Pixel = 70;
			20671: Pixel = 93;
			20672: Pixel = 119;
			20673: Pixel = 134;
			20674: Pixel = 162;
			20675: Pixel = 172;
			20676: Pixel = 151;
			20677: Pixel = 179;
			20678: Pixel = 215;
			20679: Pixel = 218;
			20680: Pixel = 193;
			20681: Pixel = 141;
			20682: Pixel = 96;
			20683: Pixel = 68;
			20684: Pixel = 63;
			20685: Pixel = 82;
			20686: Pixel = 85;
			20687: Pixel = 77;
			20688: Pixel = 84;
			20689: Pixel = 105;
			20690: Pixel = 98;
			20691: Pixel = 90;
			20692: Pixel = 93;
			20693: Pixel = 89;
			20694: Pixel = 97;
			20695: Pixel = 103;
			20696: Pixel = 95;
			20697: Pixel = 83;
			20698: Pixel = 60;
			20699: Pixel = 53;
			20700: Pixel = 45;
			20701: Pixel = 50;
			20702: Pixel = 48;
			20703: Pixel = 88;
			20704: Pixel = 160;
			20705: Pixel = 178;
			20706: Pixel = 177;
			20707: Pixel = 149;
			20708: Pixel = 71;
			20709: Pixel = 83;
			20710: Pixel = 138;
			20711: Pixel = 162;
			20712: Pixel = 172;
			20713: Pixel = 175;
			20714: Pixel = 174;
			20715: Pixel = 179;
			20716: Pixel = 178;
			20717: Pixel = 169;
			20718: Pixel = 111;
			20719: Pixel = 105;
			20720: Pixel = 83;
			20721: Pixel = 52;
			20722: Pixel = 48;
			20723: Pixel = 43;
			20724: Pixel = 43;
			20725: Pixel = 49;
			20726: Pixel = 61;
			20727: Pixel = 55;
			20728: Pixel = 48;
			20729: Pixel = 58;
			20730: Pixel = 47;
			20731: Pixel = 60;
			20732: Pixel = 63;
			20733: Pixel = 59;
			20734: Pixel = 56;
			20735: Pixel = 56;
			20736: Pixel = 50;
			20737: Pixel = 43;
			20738: Pixel = 56;
			20739: Pixel = 49;
			20740: Pixel = 47;
			20741: Pixel = 44;
			20742: Pixel = 88;
			20743: Pixel = 130;
			20744: Pixel = 137;
			20745: Pixel = 125;
			20746: Pixel = 97;
			20747: Pixel = 91;
			20748: Pixel = 90;
			20749: Pixel = 41;
			20750: Pixel = 47;
			20751: Pixel = 51;
			20752: Pixel = 44;
			20753: Pixel = 50;
			20754: Pixel = 44;
			20755: Pixel = 41;
			20756: Pixel = 39;
			20757: Pixel = 41;
			20758: Pixel = 54;
			20759: Pixel = 77;
			20760: Pixel = 99;
			20761: Pixel = 113;
			20762: Pixel = 115;
			20763: Pixel = 120;
			20764: Pixel = 113;
			20765: Pixel = 50;
			20766: Pixel = 50;
			20767: Pixel = 105;
			20768: Pixel = 129;
			20769: Pixel = 135;
			20770: Pixel = 137;
			20771: Pixel = 135;
			20772: Pixel = 138;
			20773: Pixel = 139;
			20774: Pixel = 138;
			20775: Pixel = 139;
			20776: Pixel = 142;
			20777: Pixel = 143;
			20778: Pixel = 143;
			20779: Pixel = 141;
			20780: Pixel = 140;
			20781: Pixel = 139;
			20782: Pixel = 137;
			20783: Pixel = 136;
			20784: Pixel = 136;
			20785: Pixel = 138;
			20786: Pixel = 137;
			20787: Pixel = 143;
			20788: Pixel = 144;
			20789: Pixel = 149;
			20790: Pixel = 150;
			20791: Pixel = 153;
			20792: Pixel = 155;
			20793: Pixel = 158;
			20794: Pixel = 162;
			20795: Pixel = 166;
			20796: Pixel = 174;
			20797: Pixel = 178;
			20798: Pixel = 184;
			20799: Pixel = 189;
			20800: Pixel = 196;
			20801: Pixel = 200;
			20802: Pixel = 205;
			20803: Pixel = 207;
			20804: Pixel = 209;
			20805: Pixel = 212;
			20806: Pixel = 214;
			20807: Pixel = 218;
			20808: Pixel = 211;
			20809: Pixel = 100;
			20810: Pixel = 89;
			20811: Pixel = 104;
			20812: Pixel = 100;
			20813: Pixel = 96;
			20814: Pixel = 91;
			20815: Pixel = 83;
			20816: Pixel = 72;
			20817: Pixel = 62;
			20818: Pixel = 52;
			20819: Pixel = 44;
			20820: Pixel = 41;
			20821: Pixel = 47;
			20822: Pixel = 73;
			20823: Pixel = 140;
			20824: Pixel = 198;
			20825: Pixel = 187;
			20826: Pixel = 158;
			20827: Pixel = 191;
			20828: Pixel = 215;
			20829: Pixel = 212;
			20830: Pixel = 177;
			20831: Pixel = 111;
			20832: Pixel = 71;
			20833: Pixel = 58;
			20834: Pixel = 70;
			20835: Pixel = 83;
			20836: Pixel = 72;
			20837: Pixel = 81;
			20838: Pixel = 102;
			20839: Pixel = 107;
			20840: Pixel = 93;
			20841: Pixel = 87;
			20842: Pixel = 86;
			20843: Pixel = 91;
			20844: Pixel = 101;
			20845: Pixel = 101;
			20846: Pixel = 91;
			20847: Pixel = 69;
			20848: Pixel = 55;
			20849: Pixel = 51;
			20850: Pixel = 74;
			20851: Pixel = 82;
			20852: Pixel = 75;
			20853: Pixel = 95;
			20854: Pixel = 152;
			20855: Pixel = 181;
			20856: Pixel = 183;
			20857: Pixel = 153;
			20858: Pixel = 81;
			20859: Pixel = 85;
			20860: Pixel = 135;
			20861: Pixel = 161;
			20862: Pixel = 173;
			20863: Pixel = 176;
			20864: Pixel = 174;
			20865: Pixel = 181;
			20866: Pixel = 179;
			20867: Pixel = 164;
			20868: Pixel = 111;
			20869: Pixel = 120;
			20870: Pixel = 79;
			20871: Pixel = 42;
			20872: Pixel = 48;
			20873: Pixel = 51;
			20874: Pixel = 63;
			20875: Pixel = 53;
			20876: Pixel = 43;
			20877: Pixel = 53;
			20878: Pixel = 50;
			20879: Pixel = 51;
			20880: Pixel = 57;
			20881: Pixel = 62;
			20882: Pixel = 61;
			20883: Pixel = 60;
			20884: Pixel = 60;
			20885: Pixel = 50;
			20886: Pixel = 45;
			20887: Pixel = 42;
			20888: Pixel = 45;
			20889: Pixel = 56;
			20890: Pixel = 62;
			20891: Pixel = 51;
			20892: Pixel = 38;
			20893: Pixel = 86;
			20894: Pixel = 139;
			20895: Pixel = 141;
			20896: Pixel = 104;
			20897: Pixel = 99;
			20898: Pixel = 118;
			20899: Pixel = 56;
			20900: Pixel = 46;
			20901: Pixel = 46;
			20902: Pixel = 42;
			20903: Pixel = 42;
			20904: Pixel = 42;
			20905: Pixel = 40;
			20906: Pixel = 41;
			20907: Pixel = 49;
			20908: Pixel = 73;
			20909: Pixel = 86;
			20910: Pixel = 110;
			20911: Pixel = 115;
			20912: Pixel = 119;
			20913: Pixel = 119;
			20914: Pixel = 66;
			20915: Pixel = 38;
			20916: Pixel = 86;
			20917: Pixel = 127;
			20918: Pixel = 131;
			20919: Pixel = 135;
			20920: Pixel = 134;
			20921: Pixel = 138;
			20922: Pixel = 138;
			20923: Pixel = 138;
			20924: Pixel = 139;
			20925: Pixel = 139;
			20926: Pixel = 141;
			20927: Pixel = 144;
			20928: Pixel = 143;
			20929: Pixel = 142;
			20930: Pixel = 142;
			20931: Pixel = 139;
			20932: Pixel = 137;
			20933: Pixel = 137;
			20934: Pixel = 137;
			20935: Pixel = 139;
			20936: Pixel = 138;
			20937: Pixel = 138;
			20938: Pixel = 141;
			20939: Pixel = 146;
			20940: Pixel = 146;
			20941: Pixel = 152;
			20942: Pixel = 156;
			20943: Pixel = 155;
			20944: Pixel = 159;
			20945: Pixel = 165;
			20946: Pixel = 172;
			20947: Pixel = 175;
			20948: Pixel = 182;
			20949: Pixel = 188;
			20950: Pixel = 195;
			20951: Pixel = 198;
			20952: Pixel = 203;
			20953: Pixel = 206;
			20954: Pixel = 208;
			20955: Pixel = 211;
			20956: Pixel = 213;
			20957: Pixel = 214;
			20958: Pixel = 223;
			20959: Pixel = 136;
			20960: Pixel = 82;
			20961: Pixel = 105;
			20962: Pixel = 106;
			20963: Pixel = 105;
			20964: Pixel = 99;
			20965: Pixel = 93;
			20966: Pixel = 86;
			20967: Pixel = 76;
			20968: Pixel = 61;
			20969: Pixel = 49;
			20970: Pixel = 42;
			20971: Pixel = 32;
			20972: Pixel = 63;
			20973: Pixel = 179;
			20974: Pixel = 211;
			20975: Pixel = 177;
			20976: Pixel = 159;
			20977: Pixel = 203;
			20978: Pixel = 214;
			20979: Pixel = 202;
			20980: Pixel = 137;
			20981: Pixel = 70;
			20982: Pixel = 57;
			20983: Pixel = 65;
			20984: Pixel = 78;
			20985: Pixel = 76;
			20986: Pixel = 72;
			20987: Pixel = 94;
			20988: Pixel = 110;
			20989: Pixel = 95;
			20990: Pixel = 83;
			20991: Pixel = 84;
			20992: Pixel = 82;
			20993: Pixel = 94;
			20994: Pixel = 110;
			20995: Pixel = 103;
			20996: Pixel = 85;
			20997: Pixel = 69;
			20998: Pixel = 60;
			20999: Pixel = 55;
			21000: Pixel = 92;
			21001: Pixel = 90;
			21002: Pixel = 92;
			21003: Pixel = 109;
			21004: Pixel = 150;
			21005: Pixel = 178;
			21006: Pixel = 182;
			21007: Pixel = 161;
			21008: Pixel = 96;
			21009: Pixel = 87;
			21010: Pixel = 134;
			21011: Pixel = 161;
			21012: Pixel = 173;
			21013: Pixel = 177;
			21014: Pixel = 176;
			21015: Pixel = 182;
			21016: Pixel = 181;
			21017: Pixel = 161;
			21018: Pixel = 111;
			21019: Pixel = 116;
			21020: Pixel = 85;
			21021: Pixel = 42;
			21022: Pixel = 47;
			21023: Pixel = 52;
			21024: Pixel = 53;
			21025: Pixel = 46;
			21026: Pixel = 46;
			21027: Pixel = 51;
			21028: Pixel = 53;
			21029: Pixel = 48;
			21030: Pixel = 53;
			21031: Pixel = 53;
			21032: Pixel = 63;
			21033: Pixel = 64;
			21034: Pixel = 59;
			21035: Pixel = 50;
			21036: Pixel = 44;
			21037: Pixel = 49;
			21038: Pixel = 50;
			21039: Pixel = 48;
			21040: Pixel = 68;
			21041: Pixel = 57;
			21042: Pixel = 50;
			21043: Pixel = 57;
			21044: Pixel = 84;
			21045: Pixel = 124;
			21046: Pixel = 137;
			21047: Pixel = 100;
			21048: Pixel = 100;
			21049: Pixel = 57;
			21050: Pixel = 45;
			21051: Pixel = 44;
			21052: Pixel = 43;
			21053: Pixel = 43;
			21054: Pixel = 36;
			21055: Pixel = 39;
			21056: Pixel = 45;
			21057: Pixel = 62;
			21058: Pixel = 78;
			21059: Pixel = 96;
			21060: Pixel = 116;
			21061: Pixel = 121;
			21062: Pixel = 120;
			21063: Pixel = 63;
			21064: Pixel = 37;
			21065: Pixel = 78;
			21066: Pixel = 117;
			21067: Pixel = 129;
			21068: Pixel = 132;
			21069: Pixel = 135;
			21070: Pixel = 135;
			21071: Pixel = 139;
			21072: Pixel = 140;
			21073: Pixel = 138;
			21074: Pixel = 139;
			21075: Pixel = 140;
			21076: Pixel = 140;
			21077: Pixel = 143;
			21078: Pixel = 142;
			21079: Pixel = 143;
			21080: Pixel = 143;
			21081: Pixel = 139;
			21082: Pixel = 140;
			21083: Pixel = 138;
			21084: Pixel = 136;
			21085: Pixel = 138;
			21086: Pixel = 140;
			21087: Pixel = 138;
			21088: Pixel = 140;
			21089: Pixel = 144;
			21090: Pixel = 146;
			21091: Pixel = 151;
			21092: Pixel = 153;
			21093: Pixel = 155;
			21094: Pixel = 159;
			21095: Pixel = 164;
			21096: Pixel = 167;
			21097: Pixel = 171;
			21098: Pixel = 180;
			21099: Pixel = 187;
			21100: Pixel = 192;
			21101: Pixel = 197;
			21102: Pixel = 201;
			21103: Pixel = 205;
			21104: Pixel = 207;
			21105: Pixel = 209;
			21106: Pixel = 212;
			21107: Pixel = 211;
			21108: Pixel = 223;
			21109: Pixel = 170;
			21110: Pixel = 77;
			21111: Pixel = 101;
			21112: Pixel = 108;
			21113: Pixel = 108;
			21114: Pixel = 104;
			21115: Pixel = 97;
			21116: Pixel = 91;
			21117: Pixel = 83;
			21118: Pixel = 76;
			21119: Pixel = 63;
			21120: Pixel = 49;
			21121: Pixel = 39;
			21122: Pixel = 67;
			21123: Pixel = 170;
			21124: Pixel = 205;
			21125: Pixel = 181;
			21126: Pixel = 178;
			21127: Pixel = 203;
			21128: Pixel = 201;
			21129: Pixel = 152;
			21130: Pixel = 72;
			21131: Pixel = 50;
			21132: Pixel = 59;
			21133: Pixel = 73;
			21134: Pixel = 70;
			21135: Pixel = 69;
			21136: Pixel = 89;
			21137: Pixel = 107;
			21138: Pixel = 99;
			21139: Pixel = 80;
			21140: Pixel = 77;
			21141: Pixel = 78;
			21142: Pixel = 86;
			21143: Pixel = 104;
			21144: Pixel = 113;
			21145: Pixel = 97;
			21146: Pixel = 84;
			21147: Pixel = 78;
			21148: Pixel = 61;
			21149: Pixel = 62;
			21150: Pixel = 84;
			21151: Pixel = 94;
			21152: Pixel = 104;
			21153: Pixel = 123;
			21154: Pixel = 154;
			21155: Pixel = 178;
			21156: Pixel = 181;
			21157: Pixel = 165;
			21158: Pixel = 104;
			21159: Pixel = 88;
			21160: Pixel = 132;
			21161: Pixel = 161;
			21162: Pixel = 173;
			21163: Pixel = 177;
			21164: Pixel = 177;
			21165: Pixel = 182;
			21166: Pixel = 181;
			21167: Pixel = 163;
			21168: Pixel = 105;
			21169: Pixel = 115;
			21170: Pixel = 72;
			21171: Pixel = 46;
			21172: Pixel = 49;
			21173: Pixel = 45;
			21174: Pixel = 46;
			21175: Pixel = 49;
			21176: Pixel = 46;
			21177: Pixel = 54;
			21178: Pixel = 54;
			21179: Pixel = 49;
			21180: Pixel = 46;
			21181: Pixel = 50;
			21182: Pixel = 67;
			21183: Pixel = 53;
			21184: Pixel = 61;
			21185: Pixel = 73;
			21186: Pixel = 47;
			21187: Pixel = 41;
			21188: Pixel = 69;
			21189: Pixel = 63;
			21190: Pixel = 56;
			21191: Pixel = 64;
			21192: Pixel = 57;
			21193: Pixel = 82;
			21194: Pixel = 65;
			21195: Pixel = 94;
			21196: Pixel = 89;
			21197: Pixel = 126;
			21198: Pixel = 70;
			21199: Pixel = 42;
			21200: Pixel = 47;
			21201: Pixel = 47;
			21202: Pixel = 45;
			21203: Pixel = 41;
			21204: Pixel = 38;
			21205: Pixel = 45;
			21206: Pixel = 57;
			21207: Pixel = 73;
			21208: Pixel = 90;
			21209: Pixel = 110;
			21210: Pixel = 123;
			21211: Pixel = 104;
			21212: Pixel = 54;
			21213: Pixel = 38;
			21214: Pixel = 75;
			21215: Pixel = 111;
			21216: Pixel = 125;
			21217: Pixel = 127;
			21218: Pixel = 130;
			21219: Pixel = 134;
			21220: Pixel = 136;
			21221: Pixel = 139;
			21222: Pixel = 139;
			21223: Pixel = 138;
			21224: Pixel = 138;
			21225: Pixel = 139;
			21226: Pixel = 138;
			21227: Pixel = 144;
			21228: Pixel = 142;
			21229: Pixel = 140;
			21230: Pixel = 143;
			21231: Pixel = 141;
			21232: Pixel = 141;
			21233: Pixel = 139;
			21234: Pixel = 137;
			21235: Pixel = 139;
			21236: Pixel = 141;
			21237: Pixel = 140;
			21238: Pixel = 139;
			21239: Pixel = 144;
			21240: Pixel = 145;
			21241: Pixel = 147;
			21242: Pixel = 150;
			21243: Pixel = 154;
			21244: Pixel = 159;
			21245: Pixel = 163;
			21246: Pixel = 163;
			21247: Pixel = 170;
			21248: Pixel = 175;
			21249: Pixel = 181;
			21250: Pixel = 189;
			21251: Pixel = 194;
			21252: Pixel = 199;
			21253: Pixel = 204;
			21254: Pixel = 207;
			21255: Pixel = 209;
			21256: Pixel = 212;
			21257: Pixel = 210;
			21258: Pixel = 217;
			21259: Pixel = 201;
			21260: Pixel = 92;
			21261: Pixel = 89;
			21262: Pixel = 104;
			21263: Pixel = 109;
			21264: Pixel = 105;
			21265: Pixel = 98;
			21266: Pixel = 95;
			21267: Pixel = 91;
			21268: Pixel = 83;
			21269: Pixel = 75;
			21270: Pixel = 66;
			21271: Pixel = 61;
			21272: Pixel = 75;
			21273: Pixel = 156;
			21274: Pixel = 204;
			21275: Pixel = 203;
			21276: Pixel = 193;
			21277: Pixel = 179;
			21278: Pixel = 145;
			21279: Pixel = 82;
			21280: Pixel = 51;
			21281: Pixel = 55;
			21282: Pixel = 68;
			21283: Pixel = 68;
			21284: Pixel = 66;
			21285: Pixel = 86;
			21286: Pixel = 104;
			21287: Pixel = 101;
			21288: Pixel = 87;
			21289: Pixel = 75;
			21290: Pixel = 76;
			21291: Pixel = 81;
			21292: Pixel = 99;
			21293: Pixel = 113;
			21294: Pixel = 103;
			21295: Pixel = 93;
			21296: Pixel = 83;
			21297: Pixel = 69;
			21298: Pixel = 62;
			21299: Pixel = 67;
			21300: Pixel = 71;
			21301: Pixel = 102;
			21302: Pixel = 115;
			21303: Pixel = 119;
			21304: Pixel = 149;
			21305: Pixel = 174;
			21306: Pixel = 176;
			21307: Pixel = 161;
			21308: Pixel = 108;
			21309: Pixel = 90;
			21310: Pixel = 132;
			21311: Pixel = 160;
			21312: Pixel = 173;
			21313: Pixel = 175;
			21314: Pixel = 177;
			21315: Pixel = 182;
			21316: Pixel = 179;
			21317: Pixel = 164;
			21318: Pixel = 104;
			21319: Pixel = 115;
			21320: Pixel = 65;
			21321: Pixel = 41;
			21322: Pixel = 49;
			21323: Pixel = 53;
			21324: Pixel = 50;
			21325: Pixel = 56;
			21326: Pixel = 49;
			21327: Pixel = 54;
			21328: Pixel = 57;
			21329: Pixel = 45;
			21330: Pixel = 45;
			21331: Pixel = 67;
			21332: Pixel = 84;
			21333: Pixel = 56;
			21334: Pixel = 67;
			21335: Pixel = 87;
			21336: Pixel = 48;
			21337: Pixel = 40;
			21338: Pixel = 68;
			21339: Pixel = 81;
			21340: Pixel = 54;
			21341: Pixel = 76;
			21342: Pixel = 58;
			21343: Pixel = 73;
			21344: Pixel = 73;
			21345: Pixel = 124;
			21346: Pixel = 98;
			21347: Pixel = 57;
			21348: Pixel = 81;
			21349: Pixel = 45;
			21350: Pixel = 43;
			21351: Pixel = 48;
			21352: Pixel = 41;
			21353: Pixel = 38;
			21354: Pixel = 38;
			21355: Pixel = 48;
			21356: Pixel = 73;
			21357: Pixel = 89;
			21358: Pixel = 100;
			21359: Pixel = 91;
			21360: Pixel = 66;
			21361: Pixel = 40;
			21362: Pixel = 54;
			21363: Pixel = 91;
			21364: Pixel = 111;
			21365: Pixel = 119;
			21366: Pixel = 125;
			21367: Pixel = 130;
			21368: Pixel = 132;
			21369: Pixel = 135;
			21370: Pixel = 135;
			21371: Pixel = 138;
			21372: Pixel = 137;
			21373: Pixel = 140;
			21374: Pixel = 140;
			21375: Pixel = 139;
			21376: Pixel = 141;
			21377: Pixel = 142;
			21378: Pixel = 142;
			21379: Pixel = 143;
			21380: Pixel = 144;
			21381: Pixel = 144;
			21382: Pixel = 142;
			21383: Pixel = 142;
			21384: Pixel = 140;
			21385: Pixel = 140;
			21386: Pixel = 140;
			21387: Pixel = 137;
			21388: Pixel = 138;
			21389: Pixel = 141;
			21390: Pixel = 144;
			21391: Pixel = 147;
			21392: Pixel = 148;
			21393: Pixel = 153;
			21394: Pixel = 157;
			21395: Pixel = 161;
			21396: Pixel = 165;
			21397: Pixel = 168;
			21398: Pixel = 170;
			21399: Pixel = 177;
			21400: Pixel = 185;
			21401: Pixel = 190;
			21402: Pixel = 196;
			21403: Pixel = 201;
			21404: Pixel = 205;
			21405: Pixel = 208;
			21406: Pixel = 211;
			21407: Pixel = 212;
			21408: Pixel = 213;
			21409: Pixel = 218;
			21410: Pixel = 116;
			21411: Pixel = 81;
			21412: Pixel = 101;
			21413: Pixel = 103;
			21414: Pixel = 104;
			21415: Pixel = 101;
			21416: Pixel = 97;
			21417: Pixel = 98;
			21418: Pixel = 91;
			21419: Pixel = 83;
			21420: Pixel = 85;
			21421: Pixel = 85;
			21422: Pixel = 92;
			21423: Pixel = 161;
			21424: Pixel = 210;
			21425: Pixel = 210;
			21426: Pixel = 174;
			21427: Pixel = 116;
			21428: Pixel = 77;
			21429: Pixel = 59;
			21430: Pixel = 58;
			21431: Pixel = 71;
			21432: Pixel = 73;
			21433: Pixel = 67;
			21434: Pixel = 83;
			21435: Pixel = 102;
			21436: Pixel = 106;
			21437: Pixel = 92;
			21438: Pixel = 74;
			21439: Pixel = 71;
			21440: Pixel = 78;
			21441: Pixel = 91;
			21442: Pixel = 111;
			21443: Pixel = 110;
			21444: Pixel = 99;
			21445: Pixel = 92;
			21446: Pixel = 77;
			21447: Pixel = 61;
			21448: Pixel = 70;
			21449: Pixel = 64;
			21450: Pixel = 55;
			21451: Pixel = 90;
			21452: Pixel = 101;
			21453: Pixel = 103;
			21454: Pixel = 138;
			21455: Pixel = 171;
			21456: Pixel = 179;
			21457: Pixel = 164;
			21458: Pixel = 111;
			21459: Pixel = 91;
			21460: Pixel = 129;
			21461: Pixel = 158;
			21462: Pixel = 173;
			21463: Pixel = 178;
			21464: Pixel = 179;
			21465: Pixel = 182;
			21466: Pixel = 178;
			21467: Pixel = 169;
			21468: Pixel = 106;
			21469: Pixel = 96;
			21470: Pixel = 58;
			21471: Pixel = 40;
			21472: Pixel = 48;
			21473: Pixel = 54;
			21474: Pixel = 50;
			21475: Pixel = 60;
			21476: Pixel = 49;
			21477: Pixel = 49;
			21478: Pixel = 68;
			21479: Pixel = 47;
			21480: Pixel = 47;
			21481: Pixel = 64;
			21482: Pixel = 90;
			21483: Pixel = 57;
			21484: Pixel = 67;
			21485: Pixel = 102;
			21486: Pixel = 75;
			21487: Pixel = 44;
			21488: Pixel = 59;
			21489: Pixel = 74;
			21490: Pixel = 39;
			21491: Pixel = 81;
			21492: Pixel = 90;
			21493: Pixel = 51;
			21494: Pixel = 74;
			21495: Pixel = 107;
			21496: Pixel = 142;
			21497: Pixel = 66;
			21498: Pixel = 58;
			21499: Pixel = 48;
			21500: Pixel = 40;
			21501: Pixel = 46;
			21502: Pixel = 43;
			21503: Pixel = 45;
			21504: Pixel = 44;
			21505: Pixel = 53;
			21506: Pixel = 65;
			21507: Pixel = 60;
			21508: Pixel = 50;
			21509: Pixel = 47;
			21510: Pixel = 57;
			21511: Pixel = 83;
			21512: Pixel = 105;
			21513: Pixel = 114;
			21514: Pixel = 122;
			21515: Pixel = 123;
			21516: Pixel = 126;
			21517: Pixel = 130;
			21518: Pixel = 130;
			21519: Pixel = 135;
			21520: Pixel = 136;
			21521: Pixel = 137;
			21522: Pixel = 136;
			21523: Pixel = 140;
			21524: Pixel = 139;
			21525: Pixel = 138;
			21526: Pixel = 142;
			21527: Pixel = 141;
			21528: Pixel = 143;
			21529: Pixel = 145;
			21530: Pixel = 146;
			21531: Pixel = 146;
			21532: Pixel = 145;
			21533: Pixel = 142;
			21534: Pixel = 142;
			21535: Pixel = 140;
			21536: Pixel = 138;
			21537: Pixel = 141;
			21538: Pixel = 140;
			21539: Pixel = 140;
			21540: Pixel = 143;
			21541: Pixel = 146;
			21542: Pixel = 148;
			21543: Pixel = 151;
			21544: Pixel = 154;
			21545: Pixel = 158;
			21546: Pixel = 162;
			21547: Pixel = 168;
			21548: Pixel = 173;
			21549: Pixel = 175;
			21550: Pixel = 182;
			21551: Pixel = 188;
			21552: Pixel = 194;
			21553: Pixel = 199;
			21554: Pixel = 204;
			21555: Pixel = 207;
			21556: Pixel = 210;
			21557: Pixel = 211;
			21558: Pixel = 212;
			21559: Pixel = 221;
			21560: Pixel = 150;
			21561: Pixel = 75;
			21562: Pixel = 96;
			21563: Pixel = 99;
			21564: Pixel = 102;
			21565: Pixel = 104;
			21566: Pixel = 100;
			21567: Pixel = 101;
			21568: Pixel = 96;
			21569: Pixel = 94;
			21570: Pixel = 101;
			21571: Pixel = 98;
			21572: Pixel = 95;
			21573: Pixel = 149;
			21574: Pixel = 193;
			21575: Pixel = 176;
			21576: Pixel = 111;
			21577: Pixel = 78;
			21578: Pixel = 74;
			21579: Pixel = 68;
			21580: Pixel = 74;
			21581: Pixel = 77;
			21582: Pixel = 71;
			21583: Pixel = 82;
			21584: Pixel = 105;
			21585: Pixel = 111;
			21586: Pixel = 92;
			21587: Pixel = 79;
			21588: Pixel = 69;
			21589: Pixel = 64;
			21590: Pixel = 86;
			21591: Pixel = 103;
			21592: Pixel = 113;
			21593: Pixel = 107;
			21594: Pixel = 101;
			21595: Pixel = 85;
			21596: Pixel = 63;
			21597: Pixel = 67;
			21598: Pixel = 69;
			21599: Pixel = 60;
			21600: Pixel = 47;
			21601: Pixel = 67;
			21602: Pixel = 87;
			21603: Pixel = 96;
			21604: Pixel = 131;
			21605: Pixel = 168;
			21606: Pixel = 176;
			21607: Pixel = 164;
			21608: Pixel = 121;
			21609: Pixel = 95;
			21610: Pixel = 127;
			21611: Pixel = 157;
			21612: Pixel = 172;
			21613: Pixel = 178;
			21614: Pixel = 180;
			21615: Pixel = 183;
			21616: Pixel = 180;
			21617: Pixel = 171;
			21618: Pixel = 115;
			21619: Pixel = 66;
			21620: Pixel = 48;
			21621: Pixel = 45;
			21622: Pixel = 47;
			21623: Pixel = 50;
			21624: Pixel = 51;
			21625: Pixel = 62;
			21626: Pixel = 54;
			21627: Pixel = 54;
			21628: Pixel = 73;
			21629: Pixel = 47;
			21630: Pixel = 51;
			21631: Pixel = 60;
			21632: Pixel = 85;
			21633: Pixel = 49;
			21634: Pixel = 68;
			21635: Pixel = 113;
			21636: Pixel = 105;
			21637: Pixel = 54;
			21638: Pixel = 50;
			21639: Pixel = 92;
			21640: Pixel = 51;
			21641: Pixel = 49;
			21642: Pixel = 98;
			21643: Pixel = 70;
			21644: Pixel = 69;
			21645: Pixel = 114;
			21646: Pixel = 124;
			21647: Pixel = 112;
			21648: Pixel = 58;
			21649: Pixel = 46;
			21650: Pixel = 44;
			21651: Pixel = 46;
			21652: Pixel = 47;
			21653: Pixel = 43;
			21654: Pixel = 42;
			21655: Pixel = 43;
			21656: Pixel = 47;
			21657: Pixel = 57;
			21658: Pixel = 71;
			21659: Pixel = 86;
			21660: Pixel = 103;
			21661: Pixel = 114;
			21662: Pixel = 119;
			21663: Pixel = 123;
			21664: Pixel = 125;
			21665: Pixel = 127;
			21666: Pixel = 127;
			21667: Pixel = 128;
			21668: Pixel = 129;
			21669: Pixel = 133;
			21670: Pixel = 133;
			21671: Pixel = 135;
			21672: Pixel = 137;
			21673: Pixel = 138;
			21674: Pixel = 136;
			21675: Pixel = 139;
			21676: Pixel = 140;
			21677: Pixel = 140;
			21678: Pixel = 143;
			21679: Pixel = 144;
			21680: Pixel = 146;
			21681: Pixel = 147;
			21682: Pixel = 145;
			21683: Pixel = 143;
			21684: Pixel = 143;
			21685: Pixel = 142;
			21686: Pixel = 139;
			21687: Pixel = 141;
			21688: Pixel = 142;
			21689: Pixel = 141;
			21690: Pixel = 142;
			21691: Pixel = 144;
			21692: Pixel = 149;
			21693: Pixel = 151;
			21694: Pixel = 155;
			21695: Pixel = 158;
			21696: Pixel = 161;
			21697: Pixel = 166;
			21698: Pixel = 172;
			21699: Pixel = 178;
			21700: Pixel = 182;
			21701: Pixel = 187;
			21702: Pixel = 191;
			21703: Pixel = 196;
			21704: Pixel = 201;
			21705: Pixel = 205;
			21706: Pixel = 209;
			21707: Pixel = 211;
			21708: Pixel = 211;
			21709: Pixel = 220;
			21710: Pixel = 183;
			21711: Pixel = 79;
			21712: Pixel = 87;
			21713: Pixel = 95;
			21714: Pixel = 100;
			21715: Pixel = 105;
			21716: Pixel = 107;
			21717: Pixel = 105;
			21718: Pixel = 100;
			21719: Pixel = 106;
			21720: Pixel = 112;
			21721: Pixel = 110;
			21722: Pixel = 105;
			21723: Pixel = 119;
			21724: Pixel = 135;
			21725: Pixel = 109;
			21726: Pixel = 80;
			21727: Pixel = 79;
			21728: Pixel = 82;
			21729: Pixel = 85;
			21730: Pixel = 81;
			21731: Pixel = 72;
			21732: Pixel = 78;
			21733: Pixel = 98;
			21734: Pixel = 108;
			21735: Pixel = 96;
			21736: Pixel = 76;
			21737: Pixel = 68;
			21738: Pixel = 62;
			21739: Pixel = 74;
			21740: Pixel = 102;
			21741: Pixel = 112;
			21742: Pixel = 118;
			21743: Pixel = 109;
			21744: Pixel = 97;
			21745: Pixel = 76;
			21746: Pixel = 64;
			21747: Pixel = 63;
			21748: Pixel = 60;
			21749: Pixel = 51;
			21750: Pixel = 54;
			21751: Pixel = 57;
			21752: Pixel = 75;
			21753: Pixel = 85;
			21754: Pixel = 121;
			21755: Pixel = 164;
			21756: Pixel = 178;
			21757: Pixel = 166;
			21758: Pixel = 127;
			21759: Pixel = 102;
			21760: Pixel = 125;
			21761: Pixel = 156;
			21762: Pixel = 173;
			21763: Pixel = 178;
			21764: Pixel = 180;
			21765: Pixel = 183;
			21766: Pixel = 178;
			21767: Pixel = 171;
			21768: Pixel = 114;
			21769: Pixel = 61;
			21770: Pixel = 54;
			21771: Pixel = 46;
			21772: Pixel = 53;
			21773: Pixel = 46;
			21774: Pixel = 51;
			21775: Pixel = 64;
			21776: Pixel = 59;
			21777: Pixel = 55;
			21778: Pixel = 78;
			21779: Pixel = 53;
			21780: Pixel = 44;
			21781: Pixel = 66;
			21782: Pixel = 82;
			21783: Pixel = 39;
			21784: Pixel = 61;
			21785: Pixel = 98;
			21786: Pixel = 116;
			21787: Pixel = 60;
			21788: Pixel = 37;
			21789: Pixel = 104;
			21790: Pixel = 89;
			21791: Pixel = 32;
			21792: Pixel = 74;
			21793: Pixel = 94;
			21794: Pixel = 58;
			21795: Pixel = 106;
			21796: Pixel = 104;
			21797: Pixel = 93;
			21798: Pixel = 83;
			21799: Pixel = 40;
			21800: Pixel = 49;
			21801: Pixel = 47;
			21802: Pixel = 40;
			21803: Pixel = 43;
			21804: Pixel = 50;
			21805: Pixel = 66;
			21806: Pixel = 82;
			21807: Pixel = 94;
			21808: Pixel = 103;
			21809: Pixel = 108;
			21810: Pixel = 116;
			21811: Pixel = 121;
			21812: Pixel = 123;
			21813: Pixel = 123;
			21814: Pixel = 125;
			21815: Pixel = 129;
			21816: Pixel = 128;
			21817: Pixel = 127;
			21818: Pixel = 127;
			21819: Pixel = 132;
			21820: Pixel = 134;
			21821: Pixel = 136;
			21822: Pixel = 136;
			21823: Pixel = 134;
			21824: Pixel = 139;
			21825: Pixel = 142;
			21826: Pixel = 140;
			21827: Pixel = 142;
			21828: Pixel = 141;
			21829: Pixel = 143;
			21830: Pixel = 145;
			21831: Pixel = 145;
			21832: Pixel = 143;
			21833: Pixel = 145;
			21834: Pixel = 144;
			21835: Pixel = 145;
			21836: Pixel = 143;
			21837: Pixel = 141;
			21838: Pixel = 141;
			21839: Pixel = 142;
			21840: Pixel = 143;
			21841: Pixel = 144;
			21842: Pixel = 148;
			21843: Pixel = 148;
			21844: Pixel = 153;
			21845: Pixel = 155;
			21846: Pixel = 159;
			21847: Pixel = 164;
			21848: Pixel = 168;
			21849: Pixel = 173;
			21850: Pixel = 179;
			21851: Pixel = 184;
			21852: Pixel = 188;
			21853: Pixel = 193;
			21854: Pixel = 198;
			21855: Pixel = 201;
			21856: Pixel = 208;
			21857: Pixel = 211;
			21858: Pixel = 210;
			21859: Pixel = 215;
			21860: Pixel = 207;
			21861: Pixel = 95;
			21862: Pixel = 77;
			21863: Pixel = 93;
			21864: Pixel = 98;
			21865: Pixel = 104;
			21866: Pixel = 110;
			21867: Pixel = 109;
			21868: Pixel = 109;
			21869: Pixel = 115;
			21870: Pixel = 117;
			21871: Pixel = 114;
			21872: Pixel = 114;
			21873: Pixel = 107;
			21874: Pixel = 103;
			21875: Pixel = 95;
			21876: Pixel = 91;
			21877: Pixel = 96;
			21878: Pixel = 99;
			21879: Pixel = 91;
			21880: Pixel = 80;
			21881: Pixel = 76;
			21882: Pixel = 89;
			21883: Pixel = 103;
			21884: Pixel = 94;
			21885: Pixel = 80;
			21886: Pixel = 76;
			21887: Pixel = 70;
			21888: Pixel = 65;
			21889: Pixel = 91;
			21890: Pixel = 111;
			21891: Pixel = 118;
			21892: Pixel = 115;
			21893: Pixel = 105;
			21894: Pixel = 88;
			21895: Pixel = 68;
			21896: Pixel = 60;
			21897: Pixel = 59;
			21898: Pixel = 56;
			21899: Pixel = 52;
			21900: Pixel = 55;
			21901: Pixel = 59;
			21902: Pixel = 62;
			21903: Pixel = 69;
			21904: Pixel = 114;
			21905: Pixel = 179;
			21906: Pixel = 197;
			21907: Pixel = 192;
			21908: Pixel = 148;
			21909: Pixel = 103;
			21910: Pixel = 128;
			21911: Pixel = 158;
			21912: Pixel = 174;
			21913: Pixel = 179;
			21914: Pixel = 181;
			21915: Pixel = 185;
			21916: Pixel = 184;
			21917: Pixel = 152;
			21918: Pixel = 73;
			21919: Pixel = 58;
			21920: Pixel = 58;
			21921: Pixel = 48;
			21922: Pixel = 49;
			21923: Pixel = 46;
			21924: Pixel = 53;
			21925: Pixel = 59;
			21926: Pixel = 54;
			21927: Pixel = 57;
			21928: Pixel = 65;
			21929: Pixel = 70;
			21930: Pixel = 35;
			21931: Pixel = 72;
			21932: Pixel = 86;
			21933: Pixel = 36;
			21934: Pixel = 63;
			21935: Pixel = 93;
			21936: Pixel = 99;
			21937: Pixel = 109;
			21938: Pixel = 36;
			21939: Pixel = 83;
			21940: Pixel = 113;
			21941: Pixel = 45;
			21942: Pixel = 42;
			21943: Pixel = 103;
			21944: Pixel = 72;
			21945: Pixel = 58;
			21946: Pixel = 111;
			21947: Pixel = 89;
			21948: Pixel = 50;
			21949: Pixel = 45;
			21950: Pixel = 44;
			21951: Pixel = 47;
			21952: Pixel = 48;
			21953: Pixel = 50;
			21954: Pixel = 65;
			21955: Pixel = 86;
			21956: Pixel = 99;
			21957: Pixel = 110;
			21958: Pixel = 116;
			21959: Pixel = 114;
			21960: Pixel = 118;
			21961: Pixel = 123;
			21962: Pixel = 124;
			21963: Pixel = 126;
			21964: Pixel = 128;
			21965: Pixel = 128;
			21966: Pixel = 128;
			21967: Pixel = 129;
			21968: Pixel = 129;
			21969: Pixel = 133;
			21970: Pixel = 134;
			21971: Pixel = 136;
			21972: Pixel = 135;
			21973: Pixel = 136;
			21974: Pixel = 138;
			21975: Pixel = 138;
			21976: Pixel = 138;
			21977: Pixel = 141;
			21978: Pixel = 141;
			21979: Pixel = 142;
			21980: Pixel = 144;
			21981: Pixel = 145;
			21982: Pixel = 145;
			21983: Pixel = 147;
			21984: Pixel = 144;
			21985: Pixel = 147;
			21986: Pixel = 146;
			21987: Pixel = 144;
			21988: Pixel = 144;
			21989: Pixel = 144;
			21990: Pixel = 146;
			21991: Pixel = 147;
			21992: Pixel = 148;
			21993: Pixel = 149;
			21994: Pixel = 151;
			21995: Pixel = 155;
			21996: Pixel = 159;
			21997: Pixel = 163;
			21998: Pixel = 167;
			21999: Pixel = 171;
			22000: Pixel = 177;
			22001: Pixel = 180;
			22002: Pixel = 185;
			22003: Pixel = 190;
			22004: Pixel = 197;
			22005: Pixel = 200;
			22006: Pixel = 205;
			22007: Pixel = 209;
			22008: Pixel = 208;
			22009: Pixel = 210;
			22010: Pixel = 218;
			22011: Pixel = 119;
			22012: Pixel = 70;
			22013: Pixel = 92;
			22014: Pixel = 99;
			22015: Pixel = 105;
			22016: Pixel = 109;
			22017: Pixel = 111;
			22018: Pixel = 118;
			22019: Pixel = 119;
			22020: Pixel = 118;
			22021: Pixel = 114;
			22022: Pixel = 114;
			22023: Pixel = 110;
			22024: Pixel = 105;
			22025: Pixel = 100;
			22026: Pixel = 101;
			22027: Pixel = 112;
			22028: Pixel = 105;
			22029: Pixel = 91;
			22030: Pixel = 81;
			22031: Pixel = 90;
			22032: Pixel = 99;
			22033: Pixel = 90;
			22034: Pixel = 73;
			22035: Pixel = 69;
			22036: Pixel = 73;
			22037: Pixel = 72;
			22038: Pixel = 80;
			22039: Pixel = 105;
			22040: Pixel = 120;
			22041: Pixel = 122;
			22042: Pixel = 107;
			22043: Pixel = 94;
			22044: Pixel = 76;
			22045: Pixel = 60;
			22046: Pixel = 58;
			22047: Pixel = 55;
			22048: Pixel = 51;
			22049: Pixel = 52;
			22050: Pixel = 51;
			22051: Pixel = 53;
			22052: Pixel = 56;
			22053: Pixel = 61;
			22054: Pixel = 122;
			22055: Pixel = 195;
			22056: Pixel = 204;
			22057: Pixel = 203;
			22058: Pixel = 176;
			22059: Pixel = 112;
			22060: Pixel = 126;
			22061: Pixel = 156;
			22062: Pixel = 173;
			22063: Pixel = 177;
			22064: Pixel = 179;
			22065: Pixel = 181;
			22066: Pixel = 181;
			22067: Pixel = 155;
			22068: Pixel = 101;
			22069: Pixel = 56;
			22070: Pixel = 50;
			22071: Pixel = 55;
			22072: Pixel = 49;
			22073: Pixel = 49;
			22074: Pixel = 58;
			22075: Pixel = 56;
			22076: Pixel = 58;
			22077: Pixel = 65;
			22078: Pixel = 53;
			22079: Pixel = 77;
			22080: Pixel = 39;
			22081: Pixel = 88;
			22082: Pixel = 94;
			22083: Pixel = 37;
			22084: Pixel = 69;
			22085: Pixel = 103;
			22086: Pixel = 76;
			22087: Pixel = 137;
			22088: Pixel = 60;
			22089: Pixel = 43;
			22090: Pixel = 95;
			22091: Pixel = 66;
			22092: Pixel = 45;
			22093: Pixel = 72;
			22094: Pixel = 98;
			22095: Pixel = 52;
			22096: Pixel = 79;
			22097: Pixel = 102;
			22098: Pixel = 84;
			22099: Pixel = 51;
			22100: Pixel = 32;
			22101: Pixel = 43;
			22102: Pixel = 50;
			22103: Pixel = 65;
			22104: Pixel = 85;
			22105: Pixel = 100;
			22106: Pixel = 108;
			22107: Pixel = 112;
			22108: Pixel = 117;
			22109: Pixel = 117;
			22110: Pixel = 117;
			22111: Pixel = 123;
			22112: Pixel = 126;
			22113: Pixel = 125;
			22114: Pixel = 126;
			22115: Pixel = 126;
			22116: Pixel = 129;
			22117: Pixel = 132;
			22118: Pixel = 131;
			22119: Pixel = 130;
			22120: Pixel = 132;
			22121: Pixel = 133;
			22122: Pixel = 136;
			22123: Pixel = 137;
			22124: Pixel = 135;
			22125: Pixel = 138;
			22126: Pixel = 139;
			22127: Pixel = 139;
			22128: Pixel = 140;
			22129: Pixel = 141;
			22130: Pixel = 144;
			22131: Pixel = 144;
			22132: Pixel = 146;
			22133: Pixel = 147;
			22134: Pixel = 146;
			22135: Pixel = 147;
			22136: Pixel = 147;
			22137: Pixel = 146;
			22138: Pixel = 147;
			22139: Pixel = 147;
			22140: Pixel = 146;
			22141: Pixel = 147;
			22142: Pixel = 149;
			22143: Pixel = 152;
			22144: Pixel = 151;
			22145: Pixel = 154;
			22146: Pixel = 160;
			22147: Pixel = 164;
			22148: Pixel = 167;
			22149: Pixel = 170;
			22150: Pixel = 177;
			22151: Pixel = 179;
			22152: Pixel = 185;
			22153: Pixel = 188;
			22154: Pixel = 195;
			22155: Pixel = 200;
			22156: Pixel = 203;
			22157: Pixel = 206;
			22158: Pixel = 208;
			22159: Pixel = 208;
			22160: Pixel = 221;
			22161: Pixel = 153;
			22162: Pixel = 68;
			22163: Pixel = 89;
			22164: Pixel = 97;
			22165: Pixel = 102;
			22166: Pixel = 105;
			22167: Pixel = 113;
			22168: Pixel = 120;
			22169: Pixel = 120;
			22170: Pixel = 118;
			22171: Pixel = 116;
			22172: Pixel = 114;
			22173: Pixel = 112;
			22174: Pixel = 108;
			22175: Pixel = 109;
			22176: Pixel = 118;
			22177: Pixel = 119;
			22178: Pixel = 105;
			22179: Pixel = 93;
			22180: Pixel = 95;
			22181: Pixel = 99;
			22182: Pixel = 94;
			22183: Pixel = 84;
			22184: Pixel = 74;
			22185: Pixel = 74;
			22186: Pixel = 73;
			22187: Pixel = 78;
			22188: Pixel = 101;
			22189: Pixel = 120;
			22190: Pixel = 124;
			22191: Pixel = 113;
			22192: Pixel = 101;
			22193: Pixel = 82;
			22194: Pixel = 63;
			22195: Pixel = 53;
			22196: Pixel = 58;
			22197: Pixel = 56;
			22198: Pixel = 56;
			22199: Pixel = 74;
			22200: Pixel = 49;
			22201: Pixel = 52;
			22202: Pixel = 55;
			22203: Pixel = 54;
			22204: Pixel = 124;
			22205: Pixel = 198;
			22206: Pixel = 199;
			22207: Pixel = 199;
			22208: Pixel = 184;
			22209: Pixel = 119;
			22210: Pixel = 125;
			22211: Pixel = 157;
			22212: Pixel = 173;
			22213: Pixel = 177;
			22214: Pixel = 178;
			22215: Pixel = 180;
			22216: Pixel = 181;
			22217: Pixel = 150;
			22218: Pixel = 101;
			22219: Pixel = 57;
			22220: Pixel = 48;
			22221: Pixel = 46;
			22222: Pixel = 52;
			22223: Pixel = 54;
			22224: Pixel = 60;
			22225: Pixel = 58;
			22226: Pixel = 66;
			22227: Pixel = 79;
			22228: Pixel = 63;
			22229: Pixel = 61;
			22230: Pixel = 59;
			22231: Pixel = 98;
			22232: Pixel = 77;
			22233: Pixel = 45;
			22234: Pixel = 78;
			22235: Pixel = 98;
			22236: Pixel = 62;
			22237: Pixel = 110;
			22238: Pixel = 101;
			22239: Pixel = 35;
			22240: Pixel = 102;
			22241: Pixel = 85;
			22242: Pixel = 49;
			22243: Pixel = 68;
			22244: Pixel = 80;
			22245: Pixel = 58;
			22246: Pixel = 62;
			22247: Pixel = 90;
			22248: Pixel = 101;
			22249: Pixel = 106;
			22250: Pixel = 43;
			22251: Pixel = 43;
			22252: Pixel = 64;
			22253: Pixel = 80;
			22254: Pixel = 91;
			22255: Pixel = 103;
			22256: Pixel = 109;
			22257: Pixel = 115;
			22258: Pixel = 117;
			22259: Pixel = 121;
			22260: Pixel = 121;
			22261: Pixel = 123;
			22262: Pixel = 127;
			22263: Pixel = 126;
			22264: Pixel = 126;
			22265: Pixel = 128;
			22266: Pixel = 130;
			22267: Pixel = 130;
			22268: Pixel = 131;
			22269: Pixel = 130;
			22270: Pixel = 133;
			22271: Pixel = 135;
			22272: Pixel = 137;
			22273: Pixel = 134;
			22274: Pixel = 134;
			22275: Pixel = 140;
			22276: Pixel = 139;
			22277: Pixel = 140;
			22278: Pixel = 139;
			22279: Pixel = 143;
			22280: Pixel = 144;
			22281: Pixel = 146;
			22282: Pixel = 145;
			22283: Pixel = 143;
			22284: Pixel = 146;
			22285: Pixel = 145;
			22286: Pixel = 148;
			22287: Pixel = 149;
			22288: Pixel = 148;
			22289: Pixel = 148;
			22290: Pixel = 146;
			22291: Pixel = 147;
			22292: Pixel = 150;
			22293: Pixel = 153;
			22294: Pixel = 153;
			22295: Pixel = 155;
			22296: Pixel = 160;
			22297: Pixel = 164;
			22298: Pixel = 163;
			22299: Pixel = 168;
			22300: Pixel = 173;
			22301: Pixel = 177;
			22302: Pixel = 185;
			22303: Pixel = 188;
			22304: Pixel = 193;
			22305: Pixel = 197;
			22306: Pixel = 202;
			22307: Pixel = 205;
			22308: Pixel = 208;
			22309: Pixel = 208;
			22310: Pixel = 216;
			22311: Pixel = 186;
			22312: Pixel = 77;
			22313: Pixel = 83;
			22314: Pixel = 93;
			22315: Pixel = 96;
			22316: Pixel = 101;
			22317: Pixel = 112;
			22318: Pixel = 116;
			22319: Pixel = 119;
			22320: Pixel = 126;
			22321: Pixel = 121;
			22322: Pixel = 116;
			22323: Pixel = 116;
			22324: Pixel = 119;
			22325: Pixel = 125;
			22326: Pixel = 128;
			22327: Pixel = 118;
			22328: Pixel = 100;
			22329: Pixel = 92;
			22330: Pixel = 96;
			22331: Pixel = 89;
			22332: Pixel = 80;
			22333: Pixel = 84;
			22334: Pixel = 86;
			22335: Pixel = 79;
			22336: Pixel = 79;
			22337: Pixel = 98;
			22338: Pixel = 121;
			22339: Pixel = 129;
			22340: Pixel = 122;
			22341: Pixel = 104;
			22342: Pixel = 85;
			22343: Pixel = 63;
			22344: Pixel = 51;
			22345: Pixel = 48;
			22346: Pixel = 54;
			22347: Pixel = 62;
			22348: Pixel = 80;
			22349: Pixel = 93;
			22350: Pixel = 47;
			22351: Pixel = 50;
			22352: Pixel = 52;
			22353: Pixel = 47;
			22354: Pixel = 110;
			22355: Pixel = 196;
			22356: Pixel = 198;
			22357: Pixel = 196;
			22358: Pixel = 179;
			22359: Pixel = 116;
			22360: Pixel = 128;
			22361: Pixel = 158;
			22362: Pixel = 171;
			22363: Pixel = 179;
			22364: Pixel = 180;
			22365: Pixel = 180;
			22366: Pixel = 183;
			22367: Pixel = 142;
			22368: Pixel = 76;
			22369: Pixel = 60;
			22370: Pixel = 45;
			22371: Pixel = 44;
			22372: Pixel = 57;
			22373: Pixel = 49;
			22374: Pixel = 60;
			22375: Pixel = 67;
			22376: Pixel = 66;
			22377: Pixel = 71;
			22378: Pixel = 72;
			22379: Pixel = 55;
			22380: Pixel = 86;
			22381: Pixel = 116;
			22382: Pixel = 60;
			22383: Pixel = 53;
			22384: Pixel = 74;
			22385: Pixel = 95;
			22386: Pixel = 58;
			22387: Pixel = 74;
			22388: Pixel = 111;
			22389: Pixel = 71;
			22390: Pixel = 100;
			22391: Pixel = 87;
			22392: Pixel = 36;
			22393: Pixel = 55;
			22394: Pixel = 76;
			22395: Pixel = 64;
			22396: Pixel = 43;
			22397: Pixel = 74;
			22398: Pixel = 70;
			22399: Pixel = 97;
			22400: Pixel = 90;
			22401: Pixel = 62;
			22402: Pixel = 83;
			22403: Pixel = 86;
			22404: Pixel = 93;
			22405: Pixel = 105;
			22406: Pixel = 111;
			22407: Pixel = 116;
			22408: Pixel = 119;
			22409: Pixel = 122;
			22410: Pixel = 123;
			22411: Pixel = 125;
			22412: Pixel = 127;
			22413: Pixel = 126;
			22414: Pixel = 127;
			22415: Pixel = 127;
			22416: Pixel = 128;
			22417: Pixel = 130;
			22418: Pixel = 132;
			22419: Pixel = 131;
			22420: Pixel = 130;
			22421: Pixel = 134;
			22422: Pixel = 138;
			22423: Pixel = 135;
			22424: Pixel = 133;
			22425: Pixel = 135;
			22426: Pixel = 137;
			22427: Pixel = 139;
			22428: Pixel = 141;
			22429: Pixel = 141;
			22430: Pixel = 145;
			22431: Pixel = 144;
			22432: Pixel = 144;
			22433: Pixel = 143;
			22434: Pixel = 146;
			22435: Pixel = 145;
			22436: Pixel = 146;
			22437: Pixel = 149;
			22438: Pixel = 149;
			22439: Pixel = 148;
			22440: Pixel = 149;
			22441: Pixel = 149;
			22442: Pixel = 150;
			22443: Pixel = 152;
			22444: Pixel = 156;
			22445: Pixel = 155;
			22446: Pixel = 158;
			22447: Pixel = 164;
			22448: Pixel = 164;
			22449: Pixel = 167;
			22450: Pixel = 170;
			22451: Pixel = 174;
			22452: Pixel = 182;
			22453: Pixel = 187;
			22454: Pixel = 192;
			22455: Pixel = 194;
			22456: Pixel = 199;
			22457: Pixel = 202;
			22458: Pixel = 206;
			22459: Pixel = 208;
			22460: Pixel = 213;
			22461: Pixel = 204;
			22462: Pixel = 113;
			22463: Pixel = 91;
			22464: Pixel = 91;
			22465: Pixel = 90;
			22466: Pixel = 99;
			22467: Pixel = 105;
			22468: Pixel = 114;
			22469: Pixel = 127;
			22470: Pixel = 133;
			22471: Pixel = 125;
			22472: Pixel = 123;
			22473: Pixel = 122;
			22474: Pixel = 132;
			22475: Pixel = 139;
			22476: Pixel = 128;
			22477: Pixel = 111;
			22478: Pixel = 92;
			22479: Pixel = 88;
			22480: Pixel = 79;
			22481: Pixel = 73;
			22482: Pixel = 81;
			22483: Pixel = 91;
			22484: Pixel = 88;
			22485: Pixel = 82;
			22486: Pixel = 88;
			22487: Pixel = 109;
			22488: Pixel = 127;
			22489: Pixel = 128;
			22490: Pixel = 119;
			22491: Pixel = 91;
			22492: Pixel = 64;
			22493: Pixel = 53;
			22494: Pixel = 45;
			22495: Pixel = 48;
			22496: Pixel = 58;
			22497: Pixel = 77;
			22498: Pixel = 97;
			22499: Pixel = 103;
		endcase
	end
endmodule