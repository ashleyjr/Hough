module InHandle(
	input wire			nReset,                                                      // Common to all
	input wire			Clk,                                                        // Common to all
	output reg	[7:0]	Pixel,
	output reg			Frame,
	output reg			Line
);

	parameter COLS = 102;
	parameter ROWS = 105;
	
	reg [7:0] col;
	reg [7:0] row;
	
	always @ (posedge Clk or negedge nReset) begin
		if(!nReset) begin   
			Frame <= 0;
	    	Line  <= 0;							
			row <= ROWS-1;
			col <= COLS-1;						// Zero on first pixel	
		end else begin
			if(col == (COLS-1)) begin			// Get ready for next column
	    		Line <= 1;
				col <= 0;
				row <= row + 1;
				if(row == (ROWS-1)) begin		// Get ready for next row
					Frame <= 1;
					row <= 0;
				end
			end else begin
				Line <= 0;
				Frame <= 0;
				col = col + 1;
			end
		end
	end

	always @ (*) begin
		case(col + (row*COLS))


			0: Pixel = 161;
			1: Pixel = 161;
			2: Pixel = 159;
			3: Pixel = 157;
			4: Pixel = 156;
			5: Pixel = 154;
			6: Pixel = 155;
			7: Pixel = 161;
			8: Pixel = 169;
			9: Pixel = 172;
			10: Pixel = 167;
			11: Pixel = 149;
			12: Pixel = 112;
			13: Pixel = 92;
			14: Pixel = 101;
			15: Pixel = 106;
			16: Pixel = 107;
			17: Pixel = 108;
			18: Pixel = 108;
			19: Pixel = 108;
			20: Pixel = 106;
			21: Pixel = 114;
			22: Pixel = 119;
			23: Pixel = 123;
			24: Pixel = 126;
			25: Pixel = 130;
			26: Pixel = 130;
			27: Pixel = 132;
			28: Pixel = 130;
			29: Pixel = 129;
			30: Pixel = 130;
			31: Pixel = 132;
			32: Pixel = 132;
			33: Pixel = 133;
			34: Pixel = 133;
			35: Pixel = 133;
			36: Pixel = 132;
			37: Pixel = 133;
			38: Pixel = 133;
			39: Pixel = 135;
			40: Pixel = 134;
			41: Pixel = 135;
			42: Pixel = 132;
			43: Pixel = 130;
			44: Pixel = 131;
			45: Pixel = 132;
			46: Pixel = 131;
			47: Pixel = 131;
			48: Pixel = 134;
			49: Pixel = 133;
			50: Pixel = 133;
			51: Pixel = 135;
			52: Pixel = 129;
			53: Pixel = 131;
			54: Pixel = 129;
			55: Pixel = 131;
			56: Pixel = 129;
			57: Pixel = 130;
			58: Pixel = 128;
			59: Pixel = 127;
			60: Pixel = 125;
			61: Pixel = 121;
			62: Pixel = 115;
			63: Pixel = 105;
			64: Pixel = 120;
			65: Pixel = 142;
			66: Pixel = 153;
			67: Pixel = 160;
			68: Pixel = 153;
			69: Pixel = 150;
			70: Pixel = 154;
			71: Pixel = 155;
			72: Pixel = 154;
			73: Pixel = 153;
			74: Pixel = 152;
			75: Pixel = 153;
			76: Pixel = 154;
			77: Pixel = 156;
			78: Pixel = 158;
			79: Pixel = 152;
			80: Pixel = 182;
			81: Pixel = 213;
			82: Pixel = 219;
			83: Pixel = 204;
			84: Pixel = 118;
			85: Pixel = 103;
			86: Pixel = 117;
			87: Pixel = 121;
			88: Pixel = 120;
			89: Pixel = 122;
			90: Pixel = 121;
			91: Pixel = 121;
			92: Pixel = 122;
			93: Pixel = 124;
			94: Pixel = 124;
			95: Pixel = 122;
			96: Pixel = 126;
			97: Pixel = 125;
			98: Pixel = 122;
			99: Pixel = 112;
			100: Pixel = 147;
			101: Pixel = 165;
			102: Pixel = 158;
			103: Pixel = 158;
			104: Pixel = 156;
			105: Pixel = 155;
			106: Pixel = 154;
			107: Pixel = 153;
			108: Pixel = 154;
			109: Pixel = 160;
			110: Pixel = 169;
			111: Pixel = 172;
			112: Pixel = 166;
			113: Pixel = 144;
			114: Pixel = 110;
			115: Pixel = 89;
			116: Pixel = 97;
			117: Pixel = 104;
			118: Pixel = 104;
			119: Pixel = 104;
			120: Pixel = 105;
			121: Pixel = 105;
			122: Pixel = 107;
			123: Pixel = 113;
			124: Pixel = 120;
			125: Pixel = 124;
			126: Pixel = 124;
			127: Pixel = 127;
			128: Pixel = 129;
			129: Pixel = 130;
			130: Pixel = 129;
			131: Pixel = 130;
			132: Pixel = 130;
			133: Pixel = 131;
			134: Pixel = 133;
			135: Pixel = 133;
			136: Pixel = 133;
			137: Pixel = 132;
			138: Pixel = 131;
			139: Pixel = 132;
			140: Pixel = 132;
			141: Pixel = 132;
			142: Pixel = 131;
			143: Pixel = 131;
			144: Pixel = 132;
			145: Pixel = 129;
			146: Pixel = 129;
			147: Pixel = 132;
			148: Pixel = 128;
			149: Pixel = 130;
			150: Pixel = 132;
			151: Pixel = 131;
			152: Pixel = 131;
			153: Pixel = 132;
			154: Pixel = 129;
			155: Pixel = 128;
			156: Pixel = 128;
			157: Pixel = 127;
			158: Pixel = 127;
			159: Pixel = 129;
			160: Pixel = 128;
			161: Pixel = 127;
			162: Pixel = 124;
			163: Pixel = 121;
			164: Pixel = 114;
			165: Pixel = 105;
			166: Pixel = 114;
			167: Pixel = 137;
			168: Pixel = 150;
			169: Pixel = 159;
			170: Pixel = 155;
			171: Pixel = 151;
			172: Pixel = 153;
			173: Pixel = 153;
			174: Pixel = 154;
			175: Pixel = 154;
			176: Pixel = 153;
			177: Pixel = 153;
			178: Pixel = 153;
			179: Pixel = 154;
			180: Pixel = 156;
			181: Pixel = 151;
			182: Pixel = 166;
			183: Pixel = 208;
			184: Pixel = 216;
			185: Pixel = 215;
			186: Pixel = 146;
			187: Pixel = 99;
			188: Pixel = 115;
			189: Pixel = 119;
			190: Pixel = 120;
			191: Pixel = 122;
			192: Pixel = 121;
			193: Pixel = 121;
			194: Pixel = 124;
			195: Pixel = 123;
			196: Pixel = 123;
			197: Pixel = 122;
			198: Pixel = 125;
			199: Pixel = 125;
			200: Pixel = 124;
			201: Pixel = 127;
			202: Pixel = 112;
			203: Pixel = 78;
			204: Pixel = 156;
			205: Pixel = 155;
			206: Pixel = 156;
			207: Pixel = 156;
			208: Pixel = 154;
			209: Pixel = 153;
			210: Pixel = 156;
			211: Pixel = 165;
			212: Pixel = 169;
			213: Pixel = 169;
			214: Pixel = 162;
			215: Pixel = 140;
			216: Pixel = 108;
			217: Pixel = 88;
			218: Pixel = 95;
			219: Pixel = 102;
			220: Pixel = 105;
			221: Pixel = 106;
			222: Pixel = 103;
			223: Pixel = 102;
			224: Pixel = 106;
			225: Pixel = 112;
			226: Pixel = 118;
			227: Pixel = 122;
			228: Pixel = 125;
			229: Pixel = 126;
			230: Pixel = 127;
			231: Pixel = 128;
			232: Pixel = 131;
			233: Pixel = 130;
			234: Pixel = 129;
			235: Pixel = 130;
			236: Pixel = 131;
			237: Pixel = 132;
			238: Pixel = 133;
			239: Pixel = 132;
			240: Pixel = 131;
			241: Pixel = 132;
			242: Pixel = 131;
			243: Pixel = 131;
			244: Pixel = 130;
			245: Pixel = 131;
			246: Pixel = 131;
			247: Pixel = 129;
			248: Pixel = 129;
			249: Pixel = 130;
			250: Pixel = 128;
			251: Pixel = 130;
			252: Pixel = 133;
			253: Pixel = 131;
			254: Pixel = 129;
			255: Pixel = 130;
			256: Pixel = 130;
			257: Pixel = 129;
			258: Pixel = 128;
			259: Pixel = 127;
			260: Pixel = 127;
			261: Pixel = 127;
			262: Pixel = 127;
			263: Pixel = 127;
			264: Pixel = 126;
			265: Pixel = 121;
			266: Pixel = 115;
			267: Pixel = 110;
			268: Pixel = 105;
			269: Pixel = 124;
			270: Pixel = 145;
			271: Pixel = 156;
			272: Pixel = 159;
			273: Pixel = 156;
			274: Pixel = 157;
			275: Pixel = 159;
			276: Pixel = 158;
			277: Pixel = 156;
			278: Pixel = 154;
			279: Pixel = 154;
			280: Pixel = 153;
			281: Pixel = 152;
			282: Pixel = 152;
			283: Pixel = 153;
			284: Pixel = 148;
			285: Pixel = 185;
			286: Pixel = 214;
			287: Pixel = 221;
			288: Pixel = 198;
			289: Pixel = 115;
			290: Pixel = 106;
			291: Pixel = 116;
			292: Pixel = 119;
			293: Pixel = 120;
			294: Pixel = 120;
			295: Pixel = 119;
			296: Pixel = 121;
			297: Pixel = 121;
			298: Pixel = 123;
			299: Pixel = 124;
			300: Pixel = 124;
			301: Pixel = 125;
			302: Pixel = 135;
			303: Pixel = 106;
			304: Pixel = 50;
			305: Pixel = 40;
			306: Pixel = 156;
			307: Pixel = 155;
			308: Pixel = 156;
			309: Pixel = 156;
			310: Pixel = 154;
			311: Pixel = 154;
			312: Pixel = 162;
			313: Pixel = 167;
			314: Pixel = 166;
			315: Pixel = 165;
			316: Pixel = 158;
			317: Pixel = 140;
			318: Pixel = 109;
			319: Pixel = 88;
			320: Pixel = 96;
			321: Pixel = 102;
			322: Pixel = 106;
			323: Pixel = 106;
			324: Pixel = 104;
			325: Pixel = 102;
			326: Pixel = 104;
			327: Pixel = 113;
			328: Pixel = 117;
			329: Pixel = 122;
			330: Pixel = 124;
			331: Pixel = 127;
			332: Pixel = 128;
			333: Pixel = 129;
			334: Pixel = 131;
			335: Pixel = 131;
			336: Pixel = 131;
			337: Pixel = 130;
			338: Pixel = 132;
			339: Pixel = 131;
			340: Pixel = 133;
			341: Pixel = 133;
			342: Pixel = 132;
			343: Pixel = 132;
			344: Pixel = 131;
			345: Pixel = 133;
			346: Pixel = 131;
			347: Pixel = 132;
			348: Pixel = 132;
			349: Pixel = 132;
			350: Pixel = 129;
			351: Pixel = 131;
			352: Pixel = 129;
			353: Pixel = 131;
			354: Pixel = 135;
			355: Pixel = 134;
			356: Pixel = 131;
			357: Pixel = 130;
			358: Pixel = 131;
			359: Pixel = 129;
			360: Pixel = 128;
			361: Pixel = 128;
			362: Pixel = 127;
			363: Pixel = 128;
			364: Pixel = 129;
			365: Pixel = 128;
			366: Pixel = 127;
			367: Pixel = 123;
			368: Pixel = 116;
			369: Pixel = 114;
			370: Pixel = 105;
			371: Pixel = 112;
			372: Pixel = 140;
			373: Pixel = 152;
			374: Pixel = 159;
			375: Pixel = 161;
			376: Pixel = 159;
			377: Pixel = 163;
			378: Pixel = 162;
			379: Pixel = 158;
			380: Pixel = 158;
			381: Pixel = 155;
			382: Pixel = 154;
			383: Pixel = 153;
			384: Pixel = 151;
			385: Pixel = 152;
			386: Pixel = 148;
			387: Pixel = 158;
			388: Pixel = 205;
			389: Pixel = 217;
			390: Pixel = 221;
			391: Pixel = 163;
			392: Pixel = 101;
			393: Pixel = 112;
			394: Pixel = 117;
			395: Pixel = 120;
			396: Pixel = 122;
			397: Pixel = 122;
			398: Pixel = 122;
			399: Pixel = 123;
			400: Pixel = 125;
			401: Pixel = 126;
			402: Pixel = 129;
			403: Pixel = 137;
			404: Pixel = 100;
			405: Pixel = 48;
			406: Pixel = 46;
			407: Pixel = 49;
			408: Pixel = 155;
			409: Pixel = 156;
			410: Pixel = 157;
			411: Pixel = 158;
			412: Pixel = 155;
			413: Pixel = 156;
			414: Pixel = 164;
			415: Pixel = 165;
			416: Pixel = 164;
			417: Pixel = 161;
			418: Pixel = 158;
			419: Pixel = 143;
			420: Pixel = 113;
			421: Pixel = 89;
			422: Pixel = 96;
			423: Pixel = 103;
			424: Pixel = 105;
			425: Pixel = 103;
			426: Pixel = 103;
			427: Pixel = 102;
			428: Pixel = 106;
			429: Pixel = 112;
			430: Pixel = 117;
			431: Pixel = 121;
			432: Pixel = 123;
			433: Pixel = 126;
			434: Pixel = 128;
			435: Pixel = 129;
			436: Pixel = 129;
			437: Pixel = 130;
			438: Pixel = 130;
			439: Pixel = 129;
			440: Pixel = 130;
			441: Pixel = 130;
			442: Pixel = 132;
			443: Pixel = 131;
			444: Pixel = 130;
			445: Pixel = 130;
			446: Pixel = 131;
			447: Pixel = 131;
			448: Pixel = 130;
			449: Pixel = 130;
			450: Pixel = 129;
			451: Pixel = 130;
			452: Pixel = 130;
			453: Pixel = 130;
			454: Pixel = 128;
			455: Pixel = 129;
			456: Pixel = 133;
			457: Pixel = 135;
			458: Pixel = 131;
			459: Pixel = 130;
			460: Pixel = 131;
			461: Pixel = 128;
			462: Pixel = 128;
			463: Pixel = 128;
			464: Pixel = 126;
			465: Pixel = 127;
			466: Pixel = 127;
			467: Pixel = 127;
			468: Pixel = 126;
			469: Pixel = 123;
			470: Pixel = 120;
			471: Pixel = 112;
			472: Pixel = 106;
			473: Pixel = 107;
			474: Pixel = 132;
			475: Pixel = 151;
			476: Pixel = 158;
			477: Pixel = 163;
			478: Pixel = 161;
			479: Pixel = 161;
			480: Pixel = 162;
			481: Pixel = 160;
			482: Pixel = 157;
			483: Pixel = 156;
			484: Pixel = 154;
			485: Pixel = 152;
			486: Pixel = 151;
			487: Pixel = 151;
			488: Pixel = 151;
			489: Pixel = 144;
			490: Pixel = 178;
			491: Pixel = 214;
			492: Pixel = 220;
			493: Pixel = 208;
			494: Pixel = 124;
			495: Pixel = 105;
			496: Pixel = 116;
			497: Pixel = 119;
			498: Pixel = 121;
			499: Pixel = 122;
			500: Pixel = 121;
			501: Pixel = 125;
			502: Pixel = 128;
			503: Pixel = 130;
			504: Pixel = 140;
			505: Pixel = 104;
			506: Pixel = 47;
			507: Pixel = 47;
			508: Pixel = 48;
			509: Pixel = 49;
			510: Pixel = 155;
			511: Pixel = 157;
			512: Pixel = 158;
			513: Pixel = 157;
			514: Pixel = 157;
			515: Pixel = 162;
			516: Pixel = 167;
			517: Pixel = 165;
			518: Pixel = 160;
			519: Pixel = 159;
			520: Pixel = 159;
			521: Pixel = 142;
			522: Pixel = 107;
			523: Pixel = 85;
			524: Pixel = 94;
			525: Pixel = 103;
			526: Pixel = 104;
			527: Pixel = 105;
			528: Pixel = 103;
			529: Pixel = 102;
			530: Pixel = 106;
			531: Pixel = 110;
			532: Pixel = 118;
			533: Pixel = 121;
			534: Pixel = 123;
			535: Pixel = 127;
			536: Pixel = 127;
			537: Pixel = 127;
			538: Pixel = 128;
			539: Pixel = 128;
			540: Pixel = 129;
			541: Pixel = 129;
			542: Pixel = 129;
			543: Pixel = 128;
			544: Pixel = 130;
			545: Pixel = 130;
			546: Pixel = 128;
			547: Pixel = 130;
			548: Pixel = 134;
			549: Pixel = 131;
			550: Pixel = 126;
			551: Pixel = 124;
			552: Pixel = 124;
			553: Pixel = 126;
			554: Pixel = 127;
			555: Pixel = 125;
			556: Pixel = 126;
			557: Pixel = 126;
			558: Pixel = 128;
			559: Pixel = 130;
			560: Pixel = 130;
			561: Pixel = 131;
			562: Pixel = 130;
			563: Pixel = 127;
			564: Pixel = 127;
			565: Pixel = 127;
			566: Pixel = 126;
			567: Pixel = 126;
			568: Pixel = 126;
			569: Pixel = 127;
			570: Pixel = 126;
			571: Pixel = 122;
			572: Pixel = 121;
			573: Pixel = 113;
			574: Pixel = 106;
			575: Pixel = 110;
			576: Pixel = 129;
			577: Pixel = 148;
			578: Pixel = 159;
			579: Pixel = 162;
			580: Pixel = 161;
			581: Pixel = 159;
			582: Pixel = 158;
			583: Pixel = 158;
			584: Pixel = 157;
			585: Pixel = 155;
			586: Pixel = 155;
			587: Pixel = 153;
			588: Pixel = 153;
			589: Pixel = 151;
			590: Pixel = 151;
			591: Pixel = 146;
			592: Pixel = 152;
			593: Pixel = 202;
			594: Pixel = 218;
			595: Pixel = 224;
			596: Pixel = 177;
			597: Pixel = 102;
			598: Pixel = 113;
			599: Pixel = 120;
			600: Pixel = 122;
			601: Pixel = 122;
			602: Pixel = 120;
			603: Pixel = 122;
			604: Pixel = 126;
			605: Pixel = 139;
			606: Pixel = 102;
			607: Pixel = 49;
			608: Pixel = 45;
			609: Pixel = 45;
			610: Pixel = 48;
			611: Pixel = 53;
			612: Pixel = 158;
			613: Pixel = 157;
			614: Pixel = 159;
			615: Pixel = 159;
			616: Pixel = 162;
			617: Pixel = 167;
			618: Pixel = 168;
			619: Pixel = 164;
			620: Pixel = 157;
			621: Pixel = 159;
			622: Pixel = 161;
			623: Pixel = 143;
			624: Pixel = 108;
			625: Pixel = 88;
			626: Pixel = 96;
			627: Pixel = 102;
			628: Pixel = 106;
			629: Pixel = 106;
			630: Pixel = 103;
			631: Pixel = 102;
			632: Pixel = 105;
			633: Pixel = 111;
			634: Pixel = 117;
			635: Pixel = 122;
			636: Pixel = 123;
			637: Pixel = 125;
			638: Pixel = 127;
			639: Pixel = 128;
			640: Pixel = 127;
			641: Pixel = 127;
			642: Pixel = 128;
			643: Pixel = 129;
			644: Pixel = 130;
			645: Pixel = 130;
			646: Pixel = 129;
			647: Pixel = 129;
			648: Pixel = 128;
			649: Pixel = 129;
			650: Pixel = 132;
			651: Pixel = 131;
			652: Pixel = 126;
			653: Pixel = 122;
			654: Pixel = 121;
			655: Pixel = 123;
			656: Pixel = 126;
			657: Pixel = 125;
			658: Pixel = 125;
			659: Pixel = 125;
			660: Pixel = 128;
			661: Pixel = 129;
			662: Pixel = 129;
			663: Pixel = 132;
			664: Pixel = 128;
			665: Pixel = 126;
			666: Pixel = 127;
			667: Pixel = 128;
			668: Pixel = 126;
			669: Pixel = 126;
			670: Pixel = 126;
			671: Pixel = 127;
			672: Pixel = 127;
			673: Pixel = 123;
			674: Pixel = 118;
			675: Pixel = 114;
			676: Pixel = 108;
			677: Pixel = 111;
			678: Pixel = 129;
			679: Pixel = 144;
			680: Pixel = 155;
			681: Pixel = 159;
			682: Pixel = 160;
			683: Pixel = 158;
			684: Pixel = 159;
			685: Pixel = 158;
			686: Pixel = 157;
			687: Pixel = 156;
			688: Pixel = 156;
			689: Pixel = 155;
			690: Pixel = 156;
			691: Pixel = 154;
			692: Pixel = 152;
			693: Pixel = 150;
			694: Pixel = 141;
			695: Pixel = 171;
			696: Pixel = 212;
			697: Pixel = 220;
			698: Pixel = 218;
			699: Pixel = 141;
			700: Pixel = 104;
			701: Pixel = 117;
			702: Pixel = 120;
			703: Pixel = 122;
			704: Pixel = 122;
			705: Pixel = 124;
			706: Pixel = 136;
			707: Pixel = 106;
			708: Pixel = 44;
			709: Pixel = 44;
			710: Pixel = 48;
			711: Pixel = 49;
			712: Pixel = 50;
			713: Pixel = 53;
			714: Pixel = 158;
			715: Pixel = 159;
			716: Pixel = 161;
			717: Pixel = 162;
			718: Pixel = 167;
			719: Pixel = 167;
			720: Pixel = 166;
			721: Pixel = 161;
			722: Pixel = 157;
			723: Pixel = 160;
			724: Pixel = 159;
			725: Pixel = 141;
			726: Pixel = 107;
			727: Pixel = 85;
			728: Pixel = 95;
			729: Pixel = 102;
			730: Pixel = 103;
			731: Pixel = 103;
			732: Pixel = 102;
			733: Pixel = 102;
			734: Pixel = 105;
			735: Pixel = 112;
			736: Pixel = 116;
			737: Pixel = 120;
			738: Pixel = 121;
			739: Pixel = 123;
			740: Pixel = 126;
			741: Pixel = 127;
			742: Pixel = 128;
			743: Pixel = 125;
			744: Pixel = 125;
			745: Pixel = 129;
			746: Pixel = 129;
			747: Pixel = 127;
			748: Pixel = 128;
			749: Pixel = 130;
			750: Pixel = 130;
			751: Pixel = 128;
			752: Pixel = 130;
			753: Pixel = 128;
			754: Pixel = 125;
			755: Pixel = 124;
			756: Pixel = 122;
			757: Pixel = 123;
			758: Pixel = 125;
			759: Pixel = 123;
			760: Pixel = 121;
			761: Pixel = 123;
			762: Pixel = 127;
			763: Pixel = 129;
			764: Pixel = 129;
			765: Pixel = 131;
			766: Pixel = 128;
			767: Pixel = 127;
			768: Pixel = 128;
			769: Pixel = 127;
			770: Pixel = 125;
			771: Pixel = 125;
			772: Pixel = 126;
			773: Pixel = 126;
			774: Pixel = 126;
			775: Pixel = 123;
			776: Pixel = 119;
			777: Pixel = 116;
			778: Pixel = 110;
			779: Pixel = 110;
			780: Pixel = 127;
			781: Pixel = 141;
			782: Pixel = 151;
			783: Pixel = 155;
			784: Pixel = 158;
			785: Pixel = 157;
			786: Pixel = 157;
			787: Pixel = 157;
			788: Pixel = 156;
			789: Pixel = 156;
			790: Pixel = 156;
			791: Pixel = 156;
			792: Pixel = 155;
			793: Pixel = 155;
			794: Pixel = 152;
			795: Pixel = 150;
			796: Pixel = 144;
			797: Pixel = 145;
			798: Pixel = 198;
			799: Pixel = 220;
			800: Pixel = 225;
			801: Pixel = 195;
			802: Pixel = 108;
			803: Pixel = 107;
			804: Pixel = 117;
			805: Pixel = 121;
			806: Pixel = 123;
			807: Pixel = 135;
			808: Pixel = 104;
			809: Pixel = 46;
			810: Pixel = 41;
			811: Pixel = 52;
			812: Pixel = 55;
			813: Pixel = 52;
			814: Pixel = 50;
			815: Pixel = 50;
			816: Pixel = 161;
			817: Pixel = 160;
			818: Pixel = 161;
			819: Pixel = 167;
			820: Pixel = 166;
			821: Pixel = 161;
			822: Pixel = 160;
			823: Pixel = 160;
			824: Pixel = 159;
			825: Pixel = 160;
			826: Pixel = 158;
			827: Pixel = 140;
			828: Pixel = 104;
			829: Pixel = 82;
			830: Pixel = 93;
			831: Pixel = 103;
			832: Pixel = 102;
			833: Pixel = 102;
			834: Pixel = 102;
			835: Pixel = 102;
			836: Pixel = 103;
			837: Pixel = 111;
			838: Pixel = 118;
			839: Pixel = 119;
			840: Pixel = 121;
			841: Pixel = 123;
			842: Pixel = 123;
			843: Pixel = 125;
			844: Pixel = 125;
			845: Pixel = 124;
			846: Pixel = 126;
			847: Pixel = 128;
			848: Pixel = 128;
			849: Pixel = 127;
			850: Pixel = 128;
			851: Pixel = 128;
			852: Pixel = 129;
			853: Pixel = 128;
			854: Pixel = 129;
			855: Pixel = 126;
			856: Pixel = 126;
			857: Pixel = 125;
			858: Pixel = 122;
			859: Pixel = 120;
			860: Pixel = 119;
			861: Pixel = 118;
			862: Pixel = 115;
			863: Pixel = 114;
			864: Pixel = 119;
			865: Pixel = 126;
			866: Pixel = 130;
			867: Pixel = 130;
			868: Pixel = 126;
			869: Pixel = 126;
			870: Pixel = 127;
			871: Pixel = 128;
			872: Pixel = 126;
			873: Pixel = 127;
			874: Pixel = 126;
			875: Pixel = 126;
			876: Pixel = 125;
			877: Pixel = 122;
			878: Pixel = 117;
			879: Pixel = 116;
			880: Pixel = 111;
			881: Pixel = 110;
			882: Pixel = 125;
			883: Pixel = 139;
			884: Pixel = 147;
			885: Pixel = 152;
			886: Pixel = 155;
			887: Pixel = 157;
			888: Pixel = 155;
			889: Pixel = 155;
			890: Pixel = 155;
			891: Pixel = 153;
			892: Pixel = 153;
			893: Pixel = 156;
			894: Pixel = 155;
			895: Pixel = 152;
			896: Pixel = 149;
			897: Pixel = 146;
			898: Pixel = 145;
			899: Pixel = 137;
			900: Pixel = 167;
			901: Pixel = 216;
			902: Pixel = 221;
			903: Pixel = 224;
			904: Pixel = 151;
			905: Pixel = 98;
			906: Pixel = 112;
			907: Pixel = 115;
			908: Pixel = 131;
			909: Pixel = 108;
			910: Pixel = 47;
			911: Pixel = 41;
			912: Pixel = 48;
			913: Pixel = 56;
			914: Pixel = 55;
			915: Pixel = 51;
			916: Pixel = 47;
			917: Pixel = 45;
			918: Pixel = 161;
			919: Pixel = 159;
			920: Pixel = 164;
			921: Pixel = 168;
			922: Pixel = 157;
			923: Pixel = 152;
			924: Pixel = 153;
			925: Pixel = 160;
			926: Pixel = 160;
			927: Pixel = 160;
			928: Pixel = 160;
			929: Pixel = 143;
			930: Pixel = 106;
			931: Pixel = 84;
			932: Pixel = 94;
			933: Pixel = 101;
			934: Pixel = 104;
			935: Pixel = 104;
			936: Pixel = 103;
			937: Pixel = 102;
			938: Pixel = 106;
			939: Pixel = 111;
			940: Pixel = 117;
			941: Pixel = 120;
			942: Pixel = 123;
			943: Pixel = 124;
			944: Pixel = 124;
			945: Pixel = 126;
			946: Pixel = 124;
			947: Pixel = 127;
			948: Pixel = 128;
			949: Pixel = 129;
			950: Pixel = 126;
			951: Pixel = 127;
			952: Pixel = 130;
			953: Pixel = 130;
			954: Pixel = 128;
			955: Pixel = 126;
			956: Pixel = 128;
			957: Pixel = 127;
			958: Pixel = 129;
			959: Pixel = 134;
			960: Pixel = 133;
			961: Pixel = 142;
			962: Pixel = 158;
			963: Pixel = 159;
			964: Pixel = 158;
			965: Pixel = 151;
			966: Pixel = 135;
			967: Pixel = 121;
			968: Pixel = 115;
			969: Pixel = 120;
			970: Pixel = 126;
			971: Pixel = 126;
			972: Pixel = 128;
			973: Pixel = 130;
			974: Pixel = 128;
			975: Pixel = 126;
			976: Pixel = 126;
			977: Pixel = 126;
			978: Pixel = 125;
			979: Pixel = 123;
			980: Pixel = 117;
			981: Pixel = 114;
			982: Pixel = 110;
			983: Pixel = 109;
			984: Pixel = 122;
			985: Pixel = 138;
			986: Pixel = 144;
			987: Pixel = 147;
			988: Pixel = 151;
			989: Pixel = 155;
			990: Pixel = 155;
			991: Pixel = 153;
			992: Pixel = 153;
			993: Pixel = 154;
			994: Pixel = 154;
			995: Pixel = 153;
			996: Pixel = 152;
			997: Pixel = 148;
			998: Pixel = 145;
			999: Pixel = 144;
			1000: Pixel = 143;
			1001: Pixel = 141;
			1002: Pixel = 143;
			1003: Pixel = 195;
			1004: Pixel = 220;
			1005: Pixel = 225;
			1006: Pixel = 201;
			1007: Pixel = 114;
			1008: Pixel = 106;
			1009: Pixel = 123;
			1010: Pixel = 105;
			1011: Pixel = 49;
			1012: Pixel = 43;
			1013: Pixel = 47;
			1014: Pixel = 53;
			1015: Pixel = 59;
			1016: Pixel = 55;
			1017: Pixel = 49;
			1018: Pixel = 45;
			1019: Pixel = 47;
			1020: Pixel = 161;
			1021: Pixel = 160;
			1022: Pixel = 168;
			1023: Pixel = 165;
			1024: Pixel = 148;
			1025: Pixel = 141;
			1026: Pixel = 147;
			1027: Pixel = 162;
			1028: Pixel = 161;
			1029: Pixel = 162;
			1030: Pixel = 160;
			1031: Pixel = 143;
			1032: Pixel = 107;
			1033: Pixel = 84;
			1034: Pixel = 92;
			1035: Pixel = 100;
			1036: Pixel = 104;
			1037: Pixel = 103;
			1038: Pixel = 103;
			1039: Pixel = 103;
			1040: Pixel = 107;
			1041: Pixel = 113;
			1042: Pixel = 118;
			1043: Pixel = 122;
			1044: Pixel = 121;
			1045: Pixel = 126;
			1046: Pixel = 125;
			1047: Pixel = 125;
			1048: Pixel = 127;
			1049: Pixel = 129;
			1050: Pixel = 128;
			1051: Pixel = 129;
			1052: Pixel = 128;
			1053: Pixel = 126;
			1054: Pixel = 127;
			1055: Pixel = 128;
			1056: Pixel = 127;
			1057: Pixel = 127;
			1058: Pixel = 136;
			1059: Pixel = 147;
			1060: Pixel = 145;
			1061: Pixel = 148;
			1062: Pixel = 162;
			1063: Pixel = 169;
			1064: Pixel = 177;
			1065: Pixel = 182;
			1066: Pixel = 181;
			1067: Pixel = 181;
			1068: Pixel = 185;
			1069: Pixel = 178;
			1070: Pixel = 157;
			1071: Pixel = 129;
			1072: Pixel = 114;
			1073: Pixel = 120;
			1074: Pixel = 128;
			1075: Pixel = 128;
			1076: Pixel = 128;
			1077: Pixel = 126;
			1078: Pixel = 125;
			1079: Pixel = 125;
			1080: Pixel = 124;
			1081: Pixel = 120;
			1082: Pixel = 118;
			1083: Pixel = 113;
			1084: Pixel = 109;
			1085: Pixel = 107;
			1086: Pixel = 123;
			1087: Pixel = 139;
			1088: Pixel = 144;
			1089: Pixel = 144;
			1090: Pixel = 147;
			1091: Pixel = 151;
			1092: Pixel = 154;
			1093: Pixel = 152;
			1094: Pixel = 152;
			1095: Pixel = 152;
			1096: Pixel = 152;
			1097: Pixel = 151;
			1098: Pixel = 148;
			1099: Pixel = 146;
			1100: Pixel = 143;
			1101: Pixel = 141;
			1102: Pixel = 141;
			1103: Pixel = 142;
			1104: Pixel = 138;
			1105: Pixel = 162;
			1106: Pixel = 212;
			1107: Pixel = 221;
			1108: Pixel = 227;
			1109: Pixel = 167;
			1110: Pixel = 113;
			1111: Pixel = 109;
			1112: Pixel = 47;
			1113: Pixel = 40;
			1114: Pixel = 45;
			1115: Pixel = 50;
			1116: Pixel = 54;
			1117: Pixel = 54;
			1118: Pixel = 51;
			1119: Pixel = 44;
			1120: Pixel = 46;
			1121: Pixel = 46;
			1122: Pixel = 159;
			1123: Pixel = 165;
			1124: Pixel = 169;
			1125: Pixel = 156;
			1126: Pixel = 136;
			1127: Pixel = 128;
			1128: Pixel = 148;
			1129: Pixel = 163;
			1130: Pixel = 163;
			1131: Pixel = 164;
			1132: Pixel = 161;
			1133: Pixel = 143;
			1134: Pixel = 104;
			1135: Pixel = 79;
			1136: Pixel = 91;
			1137: Pixel = 98;
			1138: Pixel = 101;
			1139: Pixel = 101;
			1140: Pixel = 102;
			1141: Pixel = 104;
			1142: Pixel = 107;
			1143: Pixel = 114;
			1144: Pixel = 118;
			1145: Pixel = 121;
			1146: Pixel = 122;
			1147: Pixel = 125;
			1148: Pixel = 124;
			1149: Pixel = 124;
			1150: Pixel = 127;
			1151: Pixel = 127;
			1152: Pixel = 128;
			1153: Pixel = 127;
			1154: Pixel = 124;
			1155: Pixel = 126;
			1156: Pixel = 134;
			1157: Pixel = 132;
			1158: Pixel = 126;
			1159: Pixel = 139;
			1160: Pixel = 145;
			1161: Pixel = 147;
			1162: Pixel = 144;
			1163: Pixel = 148;
			1164: Pixel = 156;
			1165: Pixel = 161;
			1166: Pixel = 168;
			1167: Pixel = 177;
			1168: Pixel = 174;
			1169: Pixel = 172;
			1170: Pixel = 179;
			1171: Pixel = 186;
			1172: Pixel = 195;
			1173: Pixel = 195;
			1174: Pixel = 161;
			1175: Pixel = 117;
			1176: Pixel = 114;
			1177: Pixel = 127;
			1178: Pixel = 127;
			1179: Pixel = 125;
			1180: Pixel = 125;
			1181: Pixel = 123;
			1182: Pixel = 121;
			1183: Pixel = 118;
			1184: Pixel = 114;
			1185: Pixel = 112;
			1186: Pixel = 109;
			1187: Pixel = 108;
			1188: Pixel = 124;
			1189: Pixel = 140;
			1190: Pixel = 145;
			1191: Pixel = 144;
			1192: Pixel = 146;
			1193: Pixel = 149;
			1194: Pixel = 152;
			1195: Pixel = 152;
			1196: Pixel = 149;
			1197: Pixel = 149;
			1198: Pixel = 147;
			1199: Pixel = 147;
			1200: Pixel = 144;
			1201: Pixel = 143;
			1202: Pixel = 141;
			1203: Pixel = 139;
			1204: Pixel = 139;
			1205: Pixel = 141;
			1206: Pixel = 140;
			1207: Pixel = 136;
			1208: Pixel = 185;
			1209: Pixel = 222;
			1210: Pixel = 225;
			1211: Pixel = 220;
			1212: Pixel = 134;
			1213: Pixel = 51;
			1214: Pixel = 40;
			1215: Pixel = 47;
			1216: Pixel = 51;
			1217: Pixel = 53;
			1218: Pixel = 53;
			1219: Pixel = 49;
			1220: Pixel = 48;
			1221: Pixel = 51;
			1222: Pixel = 46;
			1223: Pixel = 45;
			1224: Pixel = 163;
			1225: Pixel = 170;
			1226: Pixel = 164;
			1227: Pixel = 144;
			1228: Pixel = 113;
			1229: Pixel = 120;
			1230: Pixel = 153;
			1231: Pixel = 165;
			1232: Pixel = 165;
			1233: Pixel = 164;
			1234: Pixel = 161;
			1235: Pixel = 145;
			1236: Pixel = 105;
			1237: Pixel = 78;
			1238: Pixel = 88;
			1239: Pixel = 95;
			1240: Pixel = 98;
			1241: Pixel = 98;
			1242: Pixel = 99;
			1243: Pixel = 102;
			1244: Pixel = 106;
			1245: Pixel = 111;
			1246: Pixel = 116;
			1247: Pixel = 118;
			1248: Pixel = 121;
			1249: Pixel = 121;
			1250: Pixel = 122;
			1251: Pixel = 123;
			1252: Pixel = 125;
			1253: Pixel = 126;
			1254: Pixel = 126;
			1255: Pixel = 126;
			1256: Pixel = 134;
			1257: Pixel = 143;
			1258: Pixel = 140;
			1259: Pixel = 128;
			1260: Pixel = 122;
			1261: Pixel = 133;
			1262: Pixel = 134;
			1263: Pixel = 134;
			1264: Pixel = 143;
			1265: Pixel = 148;
			1266: Pixel = 151;
			1267: Pixel = 160;
			1268: Pixel = 164;
			1269: Pixel = 167;
			1270: Pixel = 174;
			1271: Pixel = 179;
			1272: Pixel = 183;
			1273: Pixel = 185;
			1274: Pixel = 188;
			1275: Pixel = 193;
			1276: Pixel = 201;
			1277: Pixel = 185;
			1278: Pixel = 133;
			1279: Pixel = 110;
			1280: Pixel = 119;
			1281: Pixel = 122;
			1282: Pixel = 121;
			1283: Pixel = 121;
			1284: Pixel = 120;
			1285: Pixel = 115;
			1286: Pixel = 113;
			1287: Pixel = 110;
			1288: Pixel = 105;
			1289: Pixel = 106;
			1290: Pixel = 122;
			1291: Pixel = 140;
			1292: Pixel = 147;
			1293: Pixel = 144;
			1294: Pixel = 145;
			1295: Pixel = 147;
			1296: Pixel = 148;
			1297: Pixel = 151;
			1298: Pixel = 150;
			1299: Pixel = 144;
			1300: Pixel = 143;
			1301: Pixel = 144;
			1302: Pixel = 145;
			1303: Pixel = 143;
			1304: Pixel = 142;
			1305: Pixel = 141;
			1306: Pixel = 140;
			1307: Pixel = 140;
			1308: Pixel = 143;
			1309: Pixel = 137;
			1310: Pixel = 150;
			1311: Pixel = 209;
			1312: Pixel = 222;
			1313: Pixel = 241;
			1314: Pixel = 122;
			1315: Pixel = 27;
			1316: Pixel = 47;
			1317: Pixel = 47;
			1318: Pixel = 53;
			1319: Pixel = 53;
			1320: Pixel = 50;
			1321: Pixel = 47;
			1322: Pixel = 53;
			1323: Pixel = 47;
			1324: Pixel = 47;
			1325: Pixel = 51;
			1326: Pixel = 170;
			1327: Pixel = 170;
			1328: Pixel = 155;
			1329: Pixel = 127;
			1330: Pixel = 86;
			1331: Pixel = 118;
			1332: Pixel = 154;
			1333: Pixel = 166;
			1334: Pixel = 165;
			1335: Pixel = 164;
			1336: Pixel = 161;
			1337: Pixel = 143;
			1338: Pixel = 105;
			1339: Pixel = 75;
			1340: Pixel = 83;
			1341: Pixel = 93;
			1342: Pixel = 95;
			1343: Pixel = 97;
			1344: Pixel = 100;
			1345: Pixel = 101;
			1346: Pixel = 104;
			1347: Pixel = 107;
			1348: Pixel = 114;
			1349: Pixel = 116;
			1350: Pixel = 117;
			1351: Pixel = 121;
			1352: Pixel = 123;
			1353: Pixel = 123;
			1354: Pixel = 124;
			1355: Pixel = 124;
			1356: Pixel = 123;
			1357: Pixel = 141;
			1358: Pixel = 116;
			1359: Pixel = 125;
			1360: Pixel = 120;
			1361: Pixel = 121;
			1362: Pixel = 122;
			1363: Pixel = 132;
			1364: Pixel = 128;
			1365: Pixel = 131;
			1366: Pixel = 136;
			1367: Pixel = 141;
			1368: Pixel = 147;
			1369: Pixel = 155;
			1370: Pixel = 160;
			1371: Pixel = 171;
			1372: Pixel = 176;
			1373: Pixel = 184;
			1374: Pixel = 184;
			1375: Pixel = 185;
			1376: Pixel = 187;
			1377: Pixel = 188;
			1378: Pixel = 193;
			1379: Pixel = 199;
			1380: Pixel = 197;
			1381: Pixel = 153;
			1382: Pixel = 106;
			1383: Pixel = 111;
			1384: Pixel = 119;
			1385: Pixel = 116;
			1386: Pixel = 117;
			1387: Pixel = 115;
			1388: Pixel = 111;
			1389: Pixel = 109;
			1390: Pixel = 104;
			1391: Pixel = 104;
			1392: Pixel = 122;
			1393: Pixel = 142;
			1394: Pixel = 149;
			1395: Pixel = 147;
			1396: Pixel = 144;
			1397: Pixel = 144;
			1398: Pixel = 144;
			1399: Pixel = 145;
			1400: Pixel = 151;
			1401: Pixel = 144;
			1402: Pixel = 140;
			1403: Pixel = 142;
			1404: Pixel = 145;
			1405: Pixel = 143;
			1406: Pixel = 143;
			1407: Pixel = 141;
			1408: Pixel = 140;
			1409: Pixel = 142;
			1410: Pixel = 144;
			1411: Pixel = 143;
			1412: Pixel = 138;
			1413: Pixel = 174;
			1414: Pixel = 235;
			1415: Pixel = 187;
			1416: Pixel = 49;
			1417: Pixel = 39;
			1418: Pixel = 46;
			1419: Pixel = 52;
			1420: Pixel = 55;
			1421: Pixel = 53;
			1422: Pixel = 43;
			1423: Pixel = 49;
			1424: Pixel = 48;
			1425: Pixel = 43;
			1426: Pixel = 52;
			1427: Pixel = 45;
			1428: Pixel = 172;
			1429: Pixel = 163;
			1430: Pixel = 144;
			1431: Pixel = 98;
			1432: Pixel = 77;
			1433: Pixel = 120;
			1434: Pixel = 151;
			1435: Pixel = 167;
			1436: Pixel = 165;
			1437: Pixel = 164;
			1438: Pixel = 158;
			1439: Pixel = 140;
			1440: Pixel = 103;
			1441: Pixel = 72;
			1442: Pixel = 85;
			1443: Pixel = 94;
			1444: Pixel = 100;
			1445: Pixel = 100;
			1446: Pixel = 99;
			1447: Pixel = 100;
			1448: Pixel = 103;
			1449: Pixel = 108;
			1450: Pixel = 113;
			1451: Pixel = 113;
			1452: Pixel = 116;
			1453: Pixel = 119;
			1454: Pixel = 119;
			1455: Pixel = 122;
			1456: Pixel = 124;
			1457: Pixel = 122;
			1458: Pixel = 130;
			1459: Pixel = 119;
			1460: Pixel = 112;
			1461: Pixel = 117;
			1462: Pixel = 119;
			1463: Pixel = 123;
			1464: Pixel = 123;
			1465: Pixel = 131;
			1466: Pixel = 130;
			1467: Pixel = 134;
			1468: Pixel = 133;
			1469: Pixel = 135;
			1470: Pixel = 140;
			1471: Pixel = 149;
			1472: Pixel = 163;
			1473: Pixel = 173;
			1474: Pixel = 174;
			1475: Pixel = 179;
			1476: Pixel = 182;
			1477: Pixel = 187;
			1478: Pixel = 191;
			1479: Pixel = 191;
			1480: Pixel = 195;
			1481: Pixel = 196;
			1482: Pixel = 195;
			1483: Pixel = 207;
			1484: Pixel = 176;
			1485: Pixel = 105;
			1486: Pixel = 91;
			1487: Pixel = 107;
			1488: Pixel = 113;
			1489: Pixel = 112;
			1490: Pixel = 109;
			1491: Pixel = 108;
			1492: Pixel = 105;
			1493: Pixel = 102;
			1494: Pixel = 121;
			1495: Pixel = 144;
			1496: Pixel = 152;
			1497: Pixel = 151;
			1498: Pixel = 147;
			1499: Pixel = 141;
			1500: Pixel = 138;
			1501: Pixel = 136;
			1502: Pixel = 144;
			1503: Pixel = 148;
			1504: Pixel = 142;
			1505: Pixel = 143;
			1506: Pixel = 146;
			1507: Pixel = 143;
			1508: Pixel = 142;
			1509: Pixel = 142;
			1510: Pixel = 143;
			1511: Pixel = 144;
			1512: Pixel = 144;
			1513: Pixel = 146;
			1514: Pixel = 145;
			1515: Pixel = 162;
			1516: Pixel = 172;
			1517: Pixel = 62;
			1518: Pixel = 38;
			1519: Pixel = 46;
			1520: Pixel = 48;
			1521: Pixel = 52;
			1522: Pixel = 52;
			1523: Pixel = 47;
			1524: Pixel = 52;
			1525: Pixel = 51;
			1526: Pixel = 44;
			1527: Pixel = 59;
			1528: Pixel = 53;
			1529: Pixel = 30;
			1530: Pixel = 168;
			1531: Pixel = 156;
			1532: Pixel = 122;
			1533: Pixel = 81;
			1534: Pixel = 83;
			1535: Pixel = 121;
			1536: Pixel = 152;
			1537: Pixel = 167;
			1538: Pixel = 167;
			1539: Pixel = 164;
			1540: Pixel = 158;
			1541: Pixel = 141;
			1542: Pixel = 101;
			1543: Pixel = 73;
			1544: Pixel = 85;
			1545: Pixel = 96;
			1546: Pixel = 99;
			1547: Pixel = 100;
			1548: Pixel = 99;
			1549: Pixel = 99;
			1550: Pixel = 102;
			1551: Pixel = 107;
			1552: Pixel = 112;
			1553: Pixel = 115;
			1554: Pixel = 115;
			1555: Pixel = 119;
			1556: Pixel = 119;
			1557: Pixel = 121;
			1558: Pixel = 122;
			1559: Pixel = 126;
			1560: Pixel = 140;
			1561: Pixel = 111;
			1562: Pixel = 111;
			1563: Pixel = 112;
			1564: Pixel = 117;
			1565: Pixel = 123;
			1566: Pixel = 126;
			1567: Pixel = 127;
			1568: Pixel = 132;
			1569: Pixel = 136;
			1570: Pixel = 135;
			1571: Pixel = 137;
			1572: Pixel = 139;
			1573: Pixel = 147;
			1574: Pixel = 154;
			1575: Pixel = 163;
			1576: Pixel = 174;
			1577: Pixel = 182;
			1578: Pixel = 184;
			1579: Pixel = 189;
			1580: Pixel = 190;
			1581: Pixel = 194;
			1582: Pixel = 197;
			1583: Pixel = 193;
			1584: Pixel = 191;
			1585: Pixel = 191;
			1586: Pixel = 206;
			1587: Pixel = 194;
			1588: Pixel = 148;
			1589: Pixel = 94;
			1590: Pixel = 104;
			1591: Pixel = 109;
			1592: Pixel = 105;
			1593: Pixel = 106;
			1594: Pixel = 103;
			1595: Pixel = 101;
			1596: Pixel = 122;
			1597: Pixel = 147;
			1598: Pixel = 154;
			1599: Pixel = 155;
			1600: Pixel = 151;
			1601: Pixel = 141;
			1602: Pixel = 126;
			1603: Pixel = 121;
			1604: Pixel = 135;
			1605: Pixel = 149;
			1606: Pixel = 145;
			1607: Pixel = 144;
			1608: Pixel = 147;
			1609: Pixel = 143;
			1610: Pixel = 142;
			1611: Pixel = 143;
			1612: Pixel = 144;
			1613: Pixel = 145;
			1614: Pixel = 146;
			1615: Pixel = 147;
			1616: Pixel = 154;
			1617: Pixel = 150;
			1618: Pixel = 60;
			1619: Pixel = 38;
			1620: Pixel = 44;
			1621: Pixel = 47;
			1622: Pixel = 55;
			1623: Pixel = 50;
			1624: Pixel = 44;
			1625: Pixel = 50;
			1626: Pixel = 55;
			1627: Pixel = 46;
			1628: Pixel = 57;
			1629: Pixel = 62;
			1630: Pixel = 34;
			1631: Pixel = 102;
			1632: Pixel = 160;
			1633: Pixel = 142;
			1634: Pixel = 96;
			1635: Pixel = 80;
			1636: Pixel = 86;
			1637: Pixel = 122;
			1638: Pixel = 152;
			1639: Pixel = 165;
			1640: Pixel = 168;
			1641: Pixel = 165;
			1642: Pixel = 159;
			1643: Pixel = 141;
			1644: Pixel = 100;
			1645: Pixel = 74;
			1646: Pixel = 86;
			1647: Pixel = 95;
			1648: Pixel = 99;
			1649: Pixel = 99;
			1650: Pixel = 99;
			1651: Pixel = 101;
			1652: Pixel = 103;
			1653: Pixel = 108;
			1654: Pixel = 113;
			1655: Pixel = 115;
			1656: Pixel = 116;
			1657: Pixel = 120;
			1658: Pixel = 121;
			1659: Pixel = 121;
			1660: Pixel = 120;
			1661: Pixel = 130;
			1662: Pixel = 120;
			1663: Pixel = 107;
			1664: Pixel = 110;
			1665: Pixel = 118;
			1666: Pixel = 117;
			1667: Pixel = 121;
			1668: Pixel = 123;
			1669: Pixel = 125;
			1670: Pixel = 126;
			1671: Pixel = 131;
			1672: Pixel = 134;
			1673: Pixel = 133;
			1674: Pixel = 139;
			1675: Pixel = 144;
			1676: Pixel = 152;
			1677: Pixel = 164;
			1678: Pixel = 180;
			1679: Pixel = 186;
			1680: Pixel = 185;
			1681: Pixel = 186;
			1682: Pixel = 191;
			1683: Pixel = 188;
			1684: Pixel = 186;
			1685: Pixel = 192;
			1686: Pixel = 200;
			1687: Pixel = 208;
			1688: Pixel = 212;
			1689: Pixel = 220;
			1690: Pixel = 241;
			1691: Pixel = 148;
			1692: Pixel = 79;
			1693: Pixel = 106;
			1694: Pixel = 101;
			1695: Pixel = 101;
			1696: Pixel = 100;
			1697: Pixel = 100;
			1698: Pixel = 121;
			1699: Pixel = 145;
			1700: Pixel = 154;
			1701: Pixel = 154;
			1702: Pixel = 153;
			1703: Pixel = 146;
			1704: Pixel = 117;
			1705: Pixel = 95;
			1706: Pixel = 115;
			1707: Pixel = 142;
			1708: Pixel = 148;
			1709: Pixel = 143;
			1710: Pixel = 146;
			1711: Pixel = 143;
			1712: Pixel = 143;
			1713: Pixel = 144;
			1714: Pixel = 144;
			1715: Pixel = 144;
			1716: Pixel = 146;
			1717: Pixel = 148;
			1718: Pixel = 158;
			1719: Pixel = 88;
			1720: Pixel = 39;
			1721: Pixel = 45;
			1722: Pixel = 47;
			1723: Pixel = 51;
			1724: Pixel = 52;
			1725: Pixel = 45;
			1726: Pixel = 48;
			1727: Pixel = 55;
			1728: Pixel = 46;
			1729: Pixel = 49;
			1730: Pixel = 74;
			1731: Pixel = 49;
			1732: Pixel = 84;
			1733: Pixel = 162;
			1734: Pixel = 151;
			1735: Pixel = 115;
			1736: Pixel = 82;
			1737: Pixel = 86;
			1738: Pixel = 88;
			1739: Pixel = 121;
			1740: Pixel = 151;
			1741: Pixel = 166;
			1742: Pixel = 167;
			1743: Pixel = 165;
			1744: Pixel = 158;
			1745: Pixel = 137;
			1746: Pixel = 102;
			1747: Pixel = 76;
			1748: Pixel = 86;
			1749: Pixel = 94;
			1750: Pixel = 98;
			1751: Pixel = 99;
			1752: Pixel = 102;
			1753: Pixel = 100;
			1754: Pixel = 102;
			1755: Pixel = 108;
			1756: Pixel = 113;
			1757: Pixel = 114;
			1758: Pixel = 116;
			1759: Pixel = 120;
			1760: Pixel = 121;
			1761: Pixel = 122;
			1762: Pixel = 126;
			1763: Pixel = 120;
			1764: Pixel = 105;
			1765: Pixel = 111;
			1766: Pixel = 116;
			1767: Pixel = 119;
			1768: Pixel = 121;
			1769: Pixel = 121;
			1770: Pixel = 117;
			1771: Pixel = 122;
			1772: Pixel = 129;
			1773: Pixel = 135;
			1774: Pixel = 135;
			1775: Pixel = 134;
			1776: Pixel = 138;
			1777: Pixel = 140;
			1778: Pixel = 152;
			1779: Pixel = 163;
			1780: Pixel = 177;
			1781: Pixel = 182;
			1782: Pixel = 190;
			1783: Pixel = 184;
			1784: Pixel = 176;
			1785: Pixel = 187;
			1786: Pixel = 201;
			1787: Pixel = 208;
			1788: Pixel = 210;
			1789: Pixel = 209;
			1790: Pixel = 209;
			1791: Pixel = 206;
			1792: Pixel = 217;
			1793: Pixel = 220;
			1794: Pixel = 107;
			1795: Pixel = 83;
			1796: Pixel = 100;
			1797: Pixel = 99;
			1798: Pixel = 97;
			1799: Pixel = 98;
			1800: Pixel = 119;
			1801: Pixel = 143;
			1802: Pixel = 154;
			1803: Pixel = 152;
			1804: Pixel = 153;
			1805: Pixel = 147;
			1806: Pixel = 121;
			1807: Pixel = 68;
			1808: Pixel = 82;
			1809: Pixel = 129;
			1810: Pixel = 146;
			1811: Pixel = 146;
			1812: Pixel = 145;
			1813: Pixel = 144;
			1814: Pixel = 143;
			1815: Pixel = 143;
			1816: Pixel = 144;
			1817: Pixel = 143;
			1818: Pixel = 145;
			1819: Pixel = 159;
			1820: Pixel = 117;
			1821: Pixel = 37;
			1822: Pixel = 40;
			1823: Pixel = 46;
			1824: Pixel = 53;
			1825: Pixel = 54;
			1826: Pixel = 48;
			1827: Pixel = 46;
			1828: Pixel = 53;
			1829: Pixel = 46;
			1830: Pixel = 51;
			1831: Pixel = 66;
			1832: Pixel = 67;
			1833: Pixel = 84;
			1834: Pixel = 146;
			1835: Pixel = 152;
			1836: Pixel = 131;
			1837: Pixel = 90;
			1838: Pixel = 86;
			1839: Pixel = 89;
			1840: Pixel = 87;
			1841: Pixel = 120;
			1842: Pixel = 151;
			1843: Pixel = 164;
			1844: Pixel = 166;
			1845: Pixel = 165;
			1846: Pixel = 158;
			1847: Pixel = 137;
			1848: Pixel = 102;
			1849: Pixel = 76;
			1850: Pixel = 87;
			1851: Pixel = 95;
			1852: Pixel = 96;
			1853: Pixel = 101;
			1854: Pixel = 102;
			1855: Pixel = 99;
			1856: Pixel = 103;
			1857: Pixel = 107;
			1858: Pixel = 111;
			1859: Pixel = 115;
			1860: Pixel = 117;
			1861: Pixel = 121;
			1862: Pixel = 120;
			1863: Pixel = 123;
			1864: Pixel = 121;
			1865: Pixel = 107;
			1866: Pixel = 109;
			1867: Pixel = 113;
			1868: Pixel = 117;
			1869: Pixel = 119;
			1870: Pixel = 117;
			1871: Pixel = 114;
			1872: Pixel = 120;
			1873: Pixel = 126;
			1874: Pixel = 131;
			1875: Pixel = 138;
			1876: Pixel = 137;
			1877: Pixel = 139;
			1878: Pixel = 143;
			1879: Pixel = 145;
			1880: Pixel = 148;
			1881: Pixel = 159;
			1882: Pixel = 175;
			1883: Pixel = 180;
			1884: Pixel = 169;
			1885: Pixel = 173;
			1886: Pixel = 195;
			1887: Pixel = 210;
			1888: Pixel = 209;
			1889: Pixel = 204;
			1890: Pixel = 204;
			1891: Pixel = 205;
			1892: Pixel = 205;
			1893: Pixel = 209;
			1894: Pixel = 210;
			1895: Pixel = 227;
			1896: Pixel = 201;
			1897: Pixel = 81;
			1898: Pixel = 83;
			1899: Pixel = 96;
			1900: Pixel = 94;
			1901: Pixel = 96;
			1902: Pixel = 119;
			1903: Pixel = 144;
			1904: Pixel = 155;
			1905: Pixel = 154;
			1906: Pixel = 152;
			1907: Pixel = 148;
			1908: Pixel = 127;
			1909: Pixel = 66;
			1910: Pixel = 51;
			1911: Pixel = 106;
			1912: Pixel = 137;
			1913: Pixel = 149;
			1914: Pixel = 144;
			1915: Pixel = 144;
			1916: Pixel = 142;
			1917: Pixel = 144;
			1918: Pixel = 144;
			1919: Pixel = 143;
			1920: Pixel = 152;
			1921: Pixel = 142;
			1922: Pixel = 58;
			1923: Pixel = 47;
			1924: Pixel = 45;
			1925: Pixel = 53;
			1926: Pixel = 55;
			1927: Pixel = 51;
			1928: Pixel = 45;
			1929: Pixel = 55;
			1930: Pixel = 49;
			1931: Pixel = 46;
			1932: Pixel = 62;
			1933: Pixel = 72;
			1934: Pixel = 87;
			1935: Pixel = 140;
			1936: Pixel = 150;
			1937: Pixel = 140;
			1938: Pixel = 102;
			1939: Pixel = 84;
			1940: Pixel = 93;
			1941: Pixel = 88;
			1942: Pixel = 86;
			1943: Pixel = 119;
			1944: Pixel = 149;
			1945: Pixel = 162;
			1946: Pixel = 167;
			1947: Pixel = 165;
			1948: Pixel = 159;
			1949: Pixel = 138;
			1950: Pixel = 101;
			1951: Pixel = 76;
			1952: Pixel = 89;
			1953: Pixel = 98;
			1954: Pixel = 98;
			1955: Pixel = 98;
			1956: Pixel = 99;
			1957: Pixel = 100;
			1958: Pixel = 103;
			1959: Pixel = 106;
			1960: Pixel = 113;
			1961: Pixel = 116;
			1962: Pixel = 117;
			1963: Pixel = 119;
			1964: Pixel = 122;
			1965: Pixel = 124;
			1966: Pixel = 113;
			1967: Pixel = 110;
			1968: Pixel = 113;
			1969: Pixel = 114;
			1970: Pixel = 118;
			1971: Pixel = 114;
			1972: Pixel = 112;
			1973: Pixel = 115;
			1974: Pixel = 128;
			1975: Pixel = 128;
			1976: Pixel = 134;
			1977: Pixel = 138;
			1978: Pixel = 142;
			1979: Pixel = 146;
			1980: Pixel = 140;
			1981: Pixel = 139;
			1982: Pixel = 146;
			1983: Pixel = 165;
			1984: Pixel = 167;
			1985: Pixel = 155;
			1986: Pixel = 180;
			1987: Pixel = 206;
			1988: Pixel = 204;
			1989: Pixel = 202;
			1990: Pixel = 205;
			1991: Pixel = 201;
			1992: Pixel = 199;
			1993: Pixel = 201;
			1994: Pixel = 206;
			1995: Pixel = 209;
			1996: Pixel = 209;
			1997: Pixel = 212;
			1998: Pixel = 229;
			1999: Pixel = 167;
			2000: Pixel = 76;
			2001: Pixel = 77;
			2002: Pixel = 88;
			2003: Pixel = 93;
			2004: Pixel = 120;
			2005: Pixel = 144;
			2006: Pixel = 155;
			2007: Pixel = 154;
			2008: Pixel = 153;
			2009: Pixel = 149;
			2010: Pixel = 128;
			2011: Pixel = 67;
			2012: Pixel = 41;
			2013: Pixel = 85;
			2014: Pixel = 125;
			2015: Pixel = 145;
			2016: Pixel = 147;
			2017: Pixel = 143;
			2018: Pixel = 142;
			2019: Pixel = 143;
			2020: Pixel = 144;
			2021: Pixel = 146;
			2022: Pixel = 158;
			2023: Pixel = 87;
			2024: Pixel = 34;
			2025: Pixel = 47;
			2026: Pixel = 52;
			2027: Pixel = 54;
			2028: Pixel = 51;
			2029: Pixel = 42;
			2030: Pixel = 53;
			2031: Pixel = 52;
			2032: Pixel = 49;
			2033: Pixel = 54;
			2034: Pixel = 60;
			2035: Pixel = 88;
			2036: Pixel = 135;
			2037: Pixel = 149;
			2038: Pixel = 142;
			2039: Pixel = 156;
			2040: Pixel = 86;
			2041: Pixel = 88;
			2042: Pixel = 92;
			2043: Pixel = 90;
			2044: Pixel = 87;
			2045: Pixel = 117;
			2046: Pixel = 148;
			2047: Pixel = 162;
			2048: Pixel = 166;
			2049: Pixel = 165;
			2050: Pixel = 159;
			2051: Pixel = 138;
			2052: Pixel = 103;
			2053: Pixel = 75;
			2054: Pixel = 85;
			2055: Pixel = 96;
			2056: Pixel = 99;
			2057: Pixel = 99;
			2058: Pixel = 99;
			2059: Pixel = 102;
			2060: Pixel = 103;
			2061: Pixel = 107;
			2062: Pixel = 113;
			2063: Pixel = 117;
			2064: Pixel = 117;
			2065: Pixel = 118;
			2066: Pixel = 124;
			2067: Pixel = 121;
			2068: Pixel = 109;
			2069: Pixel = 114;
			2070: Pixel = 110;
			2071: Pixel = 114;
			2072: Pixel = 116;
			2073: Pixel = 117;
			2074: Pixel = 119;
			2075: Pixel = 125;
			2076: Pixel = 128;
			2077: Pixel = 131;
			2078: Pixel = 138;
			2079: Pixel = 136;
			2080: Pixel = 140;
			2081: Pixel = 139;
			2082: Pixel = 134;
			2083: Pixel = 140;
			2084: Pixel = 146;
			2085: Pixel = 152;
			2086: Pixel = 153;
			2087: Pixel = 185;
			2088: Pixel = 201;
			2089: Pixel = 199;
			2090: Pixel = 202;
			2091: Pixel = 200;
			2092: Pixel = 198;
			2093: Pixel = 195;
			2094: Pixel = 201;
			2095: Pixel = 202;
			2096: Pixel = 203;
			2097: Pixel = 204;
			2098: Pixel = 207;
			2099: Pixel = 209;
			2100: Pixel = 210;
			2101: Pixel = 225;
			2102: Pixel = 195;
			2103: Pixel = 89;
			2104: Pixel = 72;
			2105: Pixel = 90;
			2106: Pixel = 118;
			2107: Pixel = 144;
			2108: Pixel = 155;
			2109: Pixel = 154;
			2110: Pixel = 153;
			2111: Pixel = 152;
			2112: Pixel = 126;
			2113: Pixel = 71;
			2114: Pixel = 41;
			2115: Pixel = 54;
			2116: Pixel = 101;
			2117: Pixel = 134;
			2118: Pixel = 147;
			2119: Pixel = 145;
			2120: Pixel = 141;
			2121: Pixel = 143;
			2122: Pixel = 145;
			2123: Pixel = 157;
			2124: Pixel = 122;
			2125: Pixel = 40;
			2126: Pixel = 39;
			2127: Pixel = 48;
			2128: Pixel = 57;
			2129: Pixel = 55;
			2130: Pixel = 47;
			2131: Pixel = 48;
			2132: Pixel = 55;
			2133: Pixel = 46;
			2134: Pixel = 54;
			2135: Pixel = 55;
			2136: Pixel = 69;
			2137: Pixel = 126;
			2138: Pixel = 150;
			2139: Pixel = 144;
			2140: Pixel = 156;
			2141: Pixel = 165;
			2142: Pixel = 87;
			2143: Pixel = 92;
			2144: Pixel = 92;
			2145: Pixel = 91;
			2146: Pixel = 90;
			2147: Pixel = 119;
			2148: Pixel = 148;
			2149: Pixel = 162;
			2150: Pixel = 165;
			2151: Pixel = 164;
			2152: Pixel = 158;
			2153: Pixel = 139;
			2154: Pixel = 104;
			2155: Pixel = 76;
			2156: Pixel = 85;
			2157: Pixel = 94;
			2158: Pixel = 96;
			2159: Pixel = 101;
			2160: Pixel = 99;
			2161: Pixel = 99;
			2162: Pixel = 101;
			2163: Pixel = 107;
			2164: Pixel = 112;
			2165: Pixel = 116;
			2166: Pixel = 118;
			2167: Pixel = 117;
			2168: Pixel = 137;
			2169: Pixel = 106;
			2170: Pixel = 103;
			2171: Pixel = 113;
			2172: Pixel = 113;
			2173: Pixel = 112;
			2174: Pixel = 112;
			2175: Pixel = 115;
			2176: Pixel = 121;
			2177: Pixel = 130;
			2178: Pixel = 133;
			2179: Pixel = 142;
			2180: Pixel = 137;
			2181: Pixel = 140;
			2182: Pixel = 140;
			2183: Pixel = 135;
			2184: Pixel = 133;
			2185: Pixel = 133;
			2186: Pixel = 133;
			2187: Pixel = 157;
			2188: Pixel = 191;
			2189: Pixel = 201;
			2190: Pixel = 191;
			2191: Pixel = 192;
			2192: Pixel = 191;
			2193: Pixel = 192;
			2194: Pixel = 198;
			2195: Pixel = 202;
			2196: Pixel = 202;
			2197: Pixel = 205;
			2198: Pixel = 206;
			2199: Pixel = 207;
			2200: Pixel = 207;
			2201: Pixel = 208;
			2202: Pixel = 208;
			2203: Pixel = 210;
			2204: Pixel = 229;
			2205: Pixel = 184;
			2206: Pixel = 60;
			2207: Pixel = 81;
			2208: Pixel = 116;
			2209: Pixel = 142;
			2210: Pixel = 154;
			2211: Pixel = 153;
			2212: Pixel = 153;
			2213: Pixel = 150;
			2214: Pixel = 126;
			2215: Pixel = 74;
			2216: Pixel = 42;
			2217: Pixel = 40;
			2218: Pixel = 66;
			2219: Pixel = 119;
			2220: Pixel = 142;
			2221: Pixel = 142;
			2222: Pixel = 136;
			2223: Pixel = 140;
			2224: Pixel = 150;
			2225: Pixel = 149;
			2226: Pixel = 61;
			2227: Pixel = 38;
			2228: Pixel = 46;
			2229: Pixel = 53;
			2230: Pixel = 54;
			2231: Pixel = 53;
			2232: Pixel = 47;
			2233: Pixel = 54;
			2234: Pixel = 47;
			2235: Pixel = 53;
			2236: Pixel = 51;
			2237: Pixel = 54;
			2238: Pixel = 118;
			2239: Pixel = 148;
			2240: Pixel = 137;
			2241: Pixel = 150;
			2242: Pixel = 166;
			2243: Pixel = 163;
			2244: Pixel = 90;
			2245: Pixel = 92;
			2246: Pixel = 92;
			2247: Pixel = 90;
			2248: Pixel = 88;
			2249: Pixel = 118;
			2250: Pixel = 149;
			2251: Pixel = 161;
			2252: Pixel = 164;
			2253: Pixel = 163;
			2254: Pixel = 161;
			2255: Pixel = 140;
			2256: Pixel = 103;
			2257: Pixel = 77;
			2258: Pixel = 85;
			2259: Pixel = 93;
			2260: Pixel = 97;
			2261: Pixel = 100;
			2262: Pixel = 101;
			2263: Pixel = 100;
			2264: Pixel = 103;
			2265: Pixel = 108;
			2266: Pixel = 113;
			2267: Pixel = 116;
			2268: Pixel = 109;
			2269: Pixel = 130;
			2270: Pixel = 151;
			2271: Pixel = 96;
			2272: Pixel = 108;
			2273: Pixel = 109;
			2274: Pixel = 112;
			2275: Pixel = 114;
			2276: Pixel = 116;
			2277: Pixel = 120;
			2278: Pixel = 124;
			2279: Pixel = 129;
			2280: Pixel = 139;
			2281: Pixel = 136;
			2282: Pixel = 131;
			2283: Pixel = 140;
			2284: Pixel = 139;
			2285: Pixel = 131;
			2286: Pixel = 116;
			2287: Pixel = 130;
			2288: Pixel = 170;
			2289: Pixel = 194;
			2290: Pixel = 186;
			2291: Pixel = 190;
			2292: Pixel = 191;
			2293: Pixel = 186;
			2294: Pixel = 190;
			2295: Pixel = 193;
			2296: Pixel = 199;
			2297: Pixel = 204;
			2298: Pixel = 204;
			2299: Pixel = 204;
			2300: Pixel = 204;
			2301: Pixel = 204;
			2302: Pixel = 203;
			2303: Pixel = 205;
			2304: Pixel = 204;
			2305: Pixel = 211;
			2306: Pixel = 214;
			2307: Pixel = 230;
			2308: Pixel = 131;
			2309: Pixel = 64;
			2310: Pixel = 112;
			2311: Pixel = 141;
			2312: Pixel = 152;
			2313: Pixel = 154;
			2314: Pixel = 154;
			2315: Pixel = 149;
			2316: Pixel = 127;
			2317: Pixel = 76;
			2318: Pixel = 45;
			2319: Pixel = 43;
			2320: Pixel = 44;
			2321: Pixel = 74;
			2322: Pixel = 117;
			2323: Pixel = 158;
			2324: Pixel = 153;
			2325: Pixel = 141;
			2326: Pixel = 153;
			2327: Pixel = 95;
			2328: Pixel = 37;
			2329: Pixel = 46;
			2330: Pixel = 51;
			2331: Pixel = 53;
			2332: Pixel = 55;
			2333: Pixel = 51;
			2334: Pixel = 52;
			2335: Pixel = 50;
			2336: Pixel = 52;
			2337: Pixel = 53;
			2338: Pixel = 39;
			2339: Pixel = 98;
			2340: Pixel = 152;
			2341: Pixel = 138;
			2342: Pixel = 144;
			2343: Pixel = 162;
			2344: Pixel = 161;
			2345: Pixel = 162;
			2346: Pixel = 92;
			2347: Pixel = 90;
			2348: Pixel = 90;
			2349: Pixel = 88;
			2350: Pixel = 84;
			2351: Pixel = 116;
			2352: Pixel = 149;
			2353: Pixel = 162;
			2354: Pixel = 164;
			2355: Pixel = 163;
			2356: Pixel = 161;
			2357: Pixel = 141;
			2358: Pixel = 105;
			2359: Pixel = 75;
			2360: Pixel = 84;
			2361: Pixel = 92;
			2362: Pixel = 94;
			2363: Pixel = 98;
			2364: Pixel = 99;
			2365: Pixel = 100;
			2366: Pixel = 105;
			2367: Pixel = 107;
			2368: Pixel = 111;
			2369: Pixel = 114;
			2370: Pixel = 100;
			2371: Pixel = 163;
			2372: Pixel = 138;
			2373: Pixel = 96;
			2374: Pixel = 106;
			2375: Pixel = 111;
			2376: Pixel = 112;
			2377: Pixel = 111;
			2378: Pixel = 118;
			2379: Pixel = 122;
			2380: Pixel = 129;
			2381: Pixel = 135;
			2382: Pixel = 138;
			2383: Pixel = 133;
			2384: Pixel = 134;
			2385: Pixel = 137;
			2386: Pixel = 124;
			2387: Pixel = 115;
			2388: Pixel = 133;
			2389: Pixel = 180;
			2390: Pixel = 190;
			2391: Pixel = 181;
			2392: Pixel = 189;
			2393: Pixel = 182;
			2394: Pixel = 179;
			2395: Pixel = 189;
			2396: Pixel = 198;
			2397: Pixel = 197;
			2398: Pixel = 196;
			2399: Pixel = 201;
			2400: Pixel = 203;
			2401: Pixel = 200;
			2402: Pixel = 201;
			2403: Pixel = 201;
			2404: Pixel = 200;
			2405: Pixel = 207;
			2406: Pixel = 208;
			2407: Pixel = 207;
			2408: Pixel = 210;
			2409: Pixel = 225;
			2410: Pixel = 210;
			2411: Pixel = 70;
			2412: Pixel = 105;
			2413: Pixel = 142;
			2414: Pixel = 151;
			2415: Pixel = 152;
			2416: Pixel = 154;
			2417: Pixel = 151;
			2418: Pixel = 127;
			2419: Pixel = 76;
			2420: Pixel = 45;
			2421: Pixel = 48;
			2422: Pixel = 26;
			2423: Pixel = 67;
			2424: Pixel = 185;
			2425: Pixel = 209;
			2426: Pixel = 201;
			2427: Pixel = 210;
			2428: Pixel = 167;
			2429: Pixel = 41;
			2430: Pixel = 45;
			2431: Pixel = 50;
			2432: Pixel = 55;
			2433: Pixel = 54;
			2434: Pixel = 55;
			2435: Pixel = 54;
			2436: Pixel = 51;
			2437: Pixel = 50;
			2438: Pixel = 55;
			2439: Pixel = 40;
			2440: Pixel = 74;
			2441: Pixel = 146;
			2442: Pixel = 143;
			2443: Pixel = 141;
			2444: Pixel = 161;
			2445: Pixel = 161;
			2446: Pixel = 158;
			2447: Pixel = 158;
			2448: Pixel = 89;
			2449: Pixel = 89;
			2450: Pixel = 90;
			2451: Pixel = 90;
			2452: Pixel = 85;
			2453: Pixel = 114;
			2454: Pixel = 147;
			2455: Pixel = 162;
			2456: Pixel = 164;
			2457: Pixel = 163;
			2458: Pixel = 160;
			2459: Pixel = 140;
			2460: Pixel = 101;
			2461: Pixel = 70;
			2462: Pixel = 81;
			2463: Pixel = 89;
			2464: Pixel = 95;
			2465: Pixel = 97;
			2466: Pixel = 96;
			2467: Pixel = 98;
			2468: Pixel = 102;
			2469: Pixel = 104;
			2470: Pixel = 109;
			2471: Pixel = 109;
			2472: Pixel = 107;
			2473: Pixel = 187;
			2474: Pixel = 126;
			2475: Pixel = 97;
			2476: Pixel = 108;
			2477: Pixel = 111;
			2478: Pixel = 115;
			2479: Pixel = 115;
			2480: Pixel = 117;
			2481: Pixel = 125;
			2482: Pixel = 131;
			2483: Pixel = 131;
			2484: Pixel = 127;
			2485: Pixel = 133;
			2486: Pixel = 136;
			2487: Pixel = 119;
			2488: Pixel = 108;
			2489: Pixel = 149;
			2490: Pixel = 181;
			2491: Pixel = 178;
			2492: Pixel = 179;
			2493: Pixel = 174;
			2494: Pixel = 175;
			2495: Pixel = 183;
			2496: Pixel = 186;
			2497: Pixel = 189;
			2498: Pixel = 194;
			2499: Pixel = 195;
			2500: Pixel = 195;
			2501: Pixel = 192;
			2502: Pixel = 194;
			2503: Pixel = 197;
			2504: Pixel = 202;
			2505: Pixel = 205;
			2506: Pixel = 203;
			2507: Pixel = 201;
			2508: Pixel = 206;
			2509: Pixel = 206;
			2510: Pixel = 205;
			2511: Pixel = 210;
			2512: Pixel = 231;
			2513: Pixel = 122;
			2514: Pixel = 87;
			2515: Pixel = 143;
			2516: Pixel = 152;
			2517: Pixel = 154;
			2518: Pixel = 154;
			2519: Pixel = 151;
			2520: Pixel = 126;
			2521: Pixel = 75;
			2522: Pixel = 42;
			2523: Pixel = 26;
			2524: Pixel = 87;
			2525: Pixel = 197;
			2526: Pixel = 203;
			2527: Pixel = 205;
			2528: Pixel = 220;
			2529: Pixel = 231;
			2530: Pixel = 219;
			2531: Pixel = 63;
			2532: Pixel = 39;
			2533: Pixel = 52;
			2534: Pixel = 55;
			2535: Pixel = 55;
			2536: Pixel = 50;
			2537: Pixel = 52;
			2538: Pixel = 49;
			2539: Pixel = 55;
			2540: Pixel = 49;
			2541: Pixel = 52;
			2542: Pixel = 132;
			2543: Pixel = 150;
			2544: Pixel = 140;
			2545: Pixel = 159;
			2546: Pixel = 163;
			2547: Pixel = 159;
			2548: Pixel = 158;
			2549: Pixel = 157;
			2550: Pixel = 90;
			2551: Pixel = 91;
			2552: Pixel = 94;
			2553: Pixel = 94;
			2554: Pixel = 88;
			2555: Pixel = 114;
			2556: Pixel = 146;
			2557: Pixel = 163;
			2558: Pixel = 167;
			2559: Pixel = 165;
			2560: Pixel = 159;
			2561: Pixel = 139;
			2562: Pixel = 99;
			2563: Pixel = 72;
			2564: Pixel = 78;
			2565: Pixel = 92;
			2566: Pixel = 98;
			2567: Pixel = 99;
			2568: Pixel = 100;
			2569: Pixel = 99;
			2570: Pixel = 102;
			2571: Pixel = 105;
			2572: Pixel = 112;
			2573: Pixel = 107;
			2574: Pixel = 128;
			2575: Pixel = 195;
			2576: Pixel = 114;
			2577: Pixel = 97;
			2578: Pixel = 106;
			2579: Pixel = 112;
			2580: Pixel = 110;
			2581: Pixel = 115;
			2582: Pixel = 122;
			2583: Pixel = 130;
			2584: Pixel = 121;
			2585: Pixel = 119;
			2586: Pixel = 126;
			2587: Pixel = 133;
			2588: Pixel = 117;
			2589: Pixel = 112;
			2590: Pixel = 158;
			2591: Pixel = 180;
			2592: Pixel = 171;
			2593: Pixel = 165;
			2594: Pixel = 171;
			2595: Pixel = 177;
			2596: Pixel = 178;
			2597: Pixel = 178;
			2598: Pixel = 191;
			2599: Pixel = 188;
			2600: Pixel = 189;
			2601: Pixel = 192;
			2602: Pixel = 188;
			2603: Pixel = 190;
			2604: Pixel = 196;
			2605: Pixel = 199;
			2606: Pixel = 199;
			2607: Pixel = 201;
			2608: Pixel = 199;
			2609: Pixel = 200;
			2610: Pixel = 205;
			2611: Pixel = 205;
			2612: Pixel = 206;
			2613: Pixel = 205;
			2614: Pixel = 220;
			2615: Pixel = 200;
			2616: Pixel = 95;
			2617: Pixel = 134;
			2618: Pixel = 156;
			2619: Pixel = 156;
			2620: Pixel = 155;
			2621: Pixel = 150;
			2622: Pixel = 126;
			2623: Pixel = 58;
			2624: Pixel = 24;
			2625: Pixel = 119;
			2626: Pixel = 204;
			2627: Pixel = 186;
			2628: Pixel = 206;
			2629: Pixel = 218;
			2630: Pixel = 214;
			2631: Pixel = 211;
			2632: Pixel = 237;
			2633: Pixel = 104;
			2634: Pixel = 31;
			2635: Pixel = 51;
			2636: Pixel = 54;
			2637: Pixel = 50;
			2638: Pixel = 48;
			2639: Pixel = 45;
			2640: Pixel = 50;
			2641: Pixel = 56;
			2642: Pixel = 46;
			2643: Pixel = 105;
			2644: Pixel = 155;
			2645: Pixel = 141;
			2646: Pixel = 153;
			2647: Pixel = 160;
			2648: Pixel = 158;
			2649: Pixel = 159;
			2650: Pixel = 158;
			2651: Pixel = 157;
			2652: Pixel = 94;
			2653: Pixel = 95;
			2654: Pixel = 97;
			2655: Pixel = 97;
			2656: Pixel = 94;
			2657: Pixel = 115;
			2658: Pixel = 146;
			2659: Pixel = 164;
			2660: Pixel = 167;
			2661: Pixel = 167;
			2662: Pixel = 161;
			2663: Pixel = 142;
			2664: Pixel = 102;
			2665: Pixel = 75;
			2666: Pixel = 83;
			2667: Pixel = 94;
			2668: Pixel = 98;
			2669: Pixel = 100;
			2670: Pixel = 101;
			2671: Pixel = 100;
			2672: Pixel = 105;
			2673: Pixel = 107;
			2674: Pixel = 114;
			2675: Pixel = 102;
			2676: Pixel = 146;
			2677: Pixel = 193;
			2678: Pixel = 107;
			2679: Pixel = 99;
			2680: Pixel = 106;
			2681: Pixel = 103;
			2682: Pixel = 112;
			2683: Pixel = 122;
			2684: Pixel = 125;
			2685: Pixel = 120;
			2686: Pixel = 118;
			2687: Pixel = 133;
			2688: Pixel = 134;
			2689: Pixel = 119;
			2690: Pixel = 113;
			2691: Pixel = 157;
			2692: Pixel = 172;
			2693: Pixel = 166;
			2694: Pixel = 162;
			2695: Pixel = 169;
			2696: Pixel = 178;
			2697: Pixel = 178;
			2698: Pixel = 179;
			2699: Pixel = 186;
			2700: Pixel = 184;
			2701: Pixel = 187;
			2702: Pixel = 180;
			2703: Pixel = 179;
			2704: Pixel = 187;
			2705: Pixel = 198;
			2706: Pixel = 197;
			2707: Pixel = 194;
			2708: Pixel = 193;
			2709: Pixel = 198;
			2710: Pixel = 201;
			2711: Pixel = 198;
			2712: Pixel = 198;
			2713: Pixel = 200;
			2714: Pixel = 203;
			2715: Pixel = 204;
			2716: Pixel = 205;
			2717: Pixel = 218;
			2718: Pixel = 170;
			2719: Pixel = 128;
			2720: Pixel = 152;
			2721: Pixel = 155;
			2722: Pixel = 155;
			2723: Pixel = 146;
			2724: Pixel = 98;
			2725: Pixel = 65;
			2726: Pixel = 151;
			2727: Pixel = 207;
			2728: Pixel = 185;
			2729: Pixel = 208;
			2730: Pixel = 216;
			2731: Pixel = 203;
			2732: Pixel = 202;
			2733: Pixel = 208;
			2734: Pixel = 236;
			2735: Pixel = 112;
			2736: Pixel = 31;
			2737: Pixel = 56;
			2738: Pixel = 51;
			2739: Pixel = 45;
			2740: Pixel = 46;
			2741: Pixel = 46;
			2742: Pixel = 53;
			2743: Pixel = 41;
			2744: Pixel = 67;
			2745: Pixel = 149;
			2746: Pixel = 148;
			2747: Pixel = 149;
			2748: Pixel = 161;
			2749: Pixel = 157;
			2750: Pixel = 157;
			2751: Pixel = 157;
			2752: Pixel = 155;
			2753: Pixel = 157;
			2754: Pixel = 98;
			2755: Pixel = 99;
			2756: Pixel = 100;
			2757: Pixel = 98;
			2758: Pixel = 93;
			2759: Pixel = 115;
			2760: Pixel = 147;
			2761: Pixel = 162;
			2762: Pixel = 167;
			2763: Pixel = 167;
			2764: Pixel = 164;
			2765: Pixel = 144;
			2766: Pixel = 103;
			2767: Pixel = 77;
			2768: Pixel = 85;
			2769: Pixel = 95;
			2770: Pixel = 100;
			2771: Pixel = 101;
			2772: Pixel = 103;
			2773: Pixel = 100;
			2774: Pixel = 104;
			2775: Pixel = 109;
			2776: Pixel = 115;
			2777: Pixel = 99;
			2778: Pixel = 167;
			2779: Pixel = 178;
			2780: Pixel = 103;
			2781: Pixel = 96;
			2782: Pixel = 103;
			2783: Pixel = 110;
			2784: Pixel = 113;
			2785: Pixel = 117;
			2786: Pixel = 117;
			2787: Pixel = 122;
			2788: Pixel = 127;
			2789: Pixel = 126;
			2790: Pixel = 119;
			2791: Pixel = 115;
			2792: Pixel = 155;
			2793: Pixel = 160;
			2794: Pixel = 151;
			2795: Pixel = 156;
			2796: Pixel = 165;
			2797: Pixel = 171;
			2798: Pixel = 179;
			2799: Pixel = 182;
			2800: Pixel = 177;
			2801: Pixel = 180;
			2802: Pixel = 183;
			2803: Pixel = 173;
			2804: Pixel = 174;
			2805: Pixel = 184;
			2806: Pixel = 188;
			2807: Pixel = 188;
			2808: Pixel = 195;
			2809: Pixel = 194;
			2810: Pixel = 198;
			2811: Pixel = 201;
			2812: Pixel = 186;
			2813: Pixel = 175;
			2814: Pixel = 197;
			2815: Pixel = 201;
			2816: Pixel = 202;
			2817: Pixel = 202;
			2818: Pixel = 199;
			2819: Pixel = 201;
			2820: Pixel = 219;
			2821: Pixel = 181;
			2822: Pixel = 145;
			2823: Pixel = 154;
			2824: Pixel = 147;
			2825: Pixel = 133;
			2826: Pixel = 138;
			2827: Pixel = 192;
			2828: Pixel = 202;
			2829: Pixel = 191;
			2830: Pixel = 213;
			2831: Pixel = 209;
			2832: Pixel = 202;
			2833: Pixel = 200;
			2834: Pixel = 206;
			2835: Pixel = 215;
			2836: Pixel = 232;
			2837: Pixel = 98;
			2838: Pixel = 35;
			2839: Pixel = 54;
			2840: Pixel = 54;
			2841: Pixel = 48;
			2842: Pixel = 46;
			2843: Pixel = 54;
			2844: Pixel = 48;
			2845: Pixel = 34;
			2846: Pixel = 120;
			2847: Pixel = 156;
			2848: Pixel = 145;
			2849: Pixel = 159;
			2850: Pixel = 160;
			2851: Pixel = 157;
			2852: Pixel = 156;
			2853: Pixel = 156;
			2854: Pixel = 155;
			2855: Pixel = 154;
			2856: Pixel = 99;
			2857: Pixel = 100;
			2858: Pixel = 99;
			2859: Pixel = 99;
			2860: Pixel = 97;
			2861: Pixel = 119;
			2862: Pixel = 147;
			2863: Pixel = 160;
			2864: Pixel = 168;
			2865: Pixel = 170;
			2866: Pixel = 167;
			2867: Pixel = 145;
			2868: Pixel = 104;
			2869: Pixel = 76;
			2870: Pixel = 86;
			2871: Pixel = 95;
			2872: Pixel = 99;
			2873: Pixel = 101;
			2874: Pixel = 101;
			2875: Pixel = 99;
			2876: Pixel = 101;
			2877: Pixel = 107;
			2878: Pixel = 111;
			2879: Pixel = 96;
			2880: Pixel = 180;
			2881: Pixel = 161;
			2882: Pixel = 111;
			2883: Pixel = 101;
			2884: Pixel = 105;
			2885: Pixel = 101;
			2886: Pixel = 105;
			2887: Pixel = 112;
			2888: Pixel = 118;
			2889: Pixel = 124;
			2890: Pixel = 119;
			2891: Pixel = 116;
			2892: Pixel = 118;
			2893: Pixel = 149;
			2894: Pixel = 156;
			2895: Pixel = 147;
			2896: Pixel = 145;
			2897: Pixel = 151;
			2898: Pixel = 168;
			2899: Pixel = 179;
			2900: Pixel = 172;
			2901: Pixel = 167;
			2902: Pixel = 179;
			2903: Pixel = 179;
			2904: Pixel = 169;
			2905: Pixel = 172;
			2906: Pixel = 181;
			2907: Pixel = 183;
			2908: Pixel = 181;
			2909: Pixel = 182;
			2910: Pixel = 184;
			2911: Pixel = 192;
			2912: Pixel = 196;
			2913: Pixel = 187;
			2914: Pixel = 177;
			2915: Pixel = 188;
			2916: Pixel = 194;
			2917: Pixel = 197;
			2918: Pixel = 197;
			2919: Pixel = 197;
			2920: Pixel = 196;
			2921: Pixel = 193;
			2922: Pixel = 196;
			2923: Pixel = 205;
			2924: Pixel = 156;
			2925: Pixel = 144;
			2926: Pixel = 154;
			2927: Pixel = 188;
			2928: Pixel = 204;
			2929: Pixel = 192;
			2930: Pixel = 198;
			2931: Pixel = 210;
			2932: Pixel = 203;
			2933: Pixel = 200;
			2934: Pixel = 202;
			2935: Pixel = 204;
			2936: Pixel = 210;
			2937: Pixel = 218;
			2938: Pixel = 221;
			2939: Pixel = 74;
			2940: Pixel = 43;
			2941: Pixel = 51;
			2942: Pixel = 50;
			2943: Pixel = 46;
			2944: Pixel = 45;
			2945: Pixel = 52;
			2946: Pixel = 44;
			2947: Pixel = 81;
			2948: Pixel = 152;
			2949: Pixel = 147;
			2950: Pixel = 153;
			2951: Pixel = 161;
			2952: Pixel = 158;
			2953: Pixel = 157;
			2954: Pixel = 156;
			2955: Pixel = 156;
			2956: Pixel = 154;
			2957: Pixel = 153;
			2958: Pixel = 100;
			2959: Pixel = 99;
			2960: Pixel = 99;
			2961: Pixel = 99;
			2962: Pixel = 98;
			2963: Pixel = 120;
			2964: Pixel = 149;
			2965: Pixel = 164;
			2966: Pixel = 170;
			2967: Pixel = 172;
			2968: Pixel = 170;
			2969: Pixel = 148;
			2970: Pixel = 104;
			2971: Pixel = 76;
			2972: Pixel = 88;
			2973: Pixel = 94;
			2974: Pixel = 98;
			2975: Pixel = 100;
			2976: Pixel = 100;
			2977: Pixel = 98;
			2978: Pixel = 101;
			2979: Pixel = 105;
			2980: Pixel = 103;
			2981: Pixel = 100;
			2982: Pixel = 194;
			2983: Pixel = 161;
			2984: Pixel = 118;
			2985: Pixel = 102;
			2986: Pixel = 105;
			2987: Pixel = 104;
			2988: Pixel = 108;
			2989: Pixel = 112;
			2990: Pixel = 117;
			2991: Pixel = 119;
			2992: Pixel = 120;
			2993: Pixel = 121;
			2994: Pixel = 152;
			2995: Pixel = 147;
			2996: Pixel = 144;
			2997: Pixel = 141;
			2998: Pixel = 146;
			2999: Pixel = 163;
			3000: Pixel = 164;
			3001: Pixel = 165;
			3002: Pixel = 169;
			3003: Pixel = 172;
			3004: Pixel = 171;
			3005: Pixel = 165;
			3006: Pixel = 169;
			3007: Pixel = 178;
			3008: Pixel = 175;
			3009: Pixel = 176;
			3010: Pixel = 176;
			3011: Pixel = 179;
			3012: Pixel = 186;
			3013: Pixel = 179;
			3014: Pixel = 174;
			3015: Pixel = 184;
			3016: Pixel = 183;
			3017: Pixel = 185;
			3018: Pixel = 190;
			3019: Pixel = 194;
			3020: Pixel = 190;
			3021: Pixel = 186;
			3022: Pixel = 190;
			3023: Pixel = 188;
			3024: Pixel = 185;
			3025: Pixel = 192;
			3026: Pixel = 174;
			3027: Pixel = 174;
			3028: Pixel = 198;
			3029: Pixel = 195;
			3030: Pixel = 193;
			3031: Pixel = 204;
			3032: Pixel = 207;
			3033: Pixel = 199;
			3034: Pixel = 200;
			3035: Pixel = 203;
			3036: Pixel = 204;
			3037: Pixel = 202;
			3038: Pixel = 207;
			3039: Pixel = 223;
			3040: Pixel = 206;
			3041: Pixel = 54;
			3042: Pixel = 48;
			3043: Pixel = 54;
			3044: Pixel = 50;
			3045: Pixel = 43;
			3046: Pixel = 49;
			3047: Pixel = 54;
			3048: Pixel = 68;
			3049: Pixel = 131;
			3050: Pixel = 150;
			3051: Pixel = 147;
			3052: Pixel = 160;
			3053: Pixel = 159;
			3054: Pixel = 158;
			3055: Pixel = 156;
			3056: Pixel = 157;
			3057: Pixel = 154;
			3058: Pixel = 154;
			3059: Pixel = 153;
			3060: Pixel = 99;
			3061: Pixel = 99;
			3062: Pixel = 98;
			3063: Pixel = 98;
			3064: Pixel = 99;
			3065: Pixel = 118;
			3066: Pixel = 148;
			3067: Pixel = 166;
			3068: Pixel = 172;
			3069: Pixel = 174;
			3070: Pixel = 170;
			3071: Pixel = 147;
			3072: Pixel = 105;
			3073: Pixel = 75;
			3074: Pixel = 84;
			3075: Pixel = 94;
			3076: Pixel = 97;
			3077: Pixel = 99;
			3078: Pixel = 98;
			3079: Pixel = 98;
			3080: Pixel = 99;
			3081: Pixel = 105;
			3082: Pixel = 98;
			3083: Pixel = 111;
			3084: Pixel = 205;
			3085: Pixel = 163;
			3086: Pixel = 128;
			3087: Pixel = 112;
			3088: Pixel = 107;
			3089: Pixel = 105;
			3090: Pixel = 111;
			3091: Pixel = 114;
			3092: Pixel = 122;
			3093: Pixel = 122;
			3094: Pixel = 117;
			3095: Pixel = 146;
			3096: Pixel = 144;
			3097: Pixel = 145;
			3098: Pixel = 135;
			3099: Pixel = 140;
			3100: Pixel = 152;
			3101: Pixel = 155;
			3102: Pixel = 155;
			3103: Pixel = 165;
			3104: Pixel = 174;
			3105: Pixel = 168;
			3106: Pixel = 160;
			3107: Pixel = 173;
			3108: Pixel = 174;
			3109: Pixel = 172;
			3110: Pixel = 175;
			3111: Pixel = 173;
			3112: Pixel = 171;
			3113: Pixel = 181;
			3114: Pixel = 184;
			3115: Pixel = 181;
			3116: Pixel = 181;
			3117: Pixel = 183;
			3118: Pixel = 188;
			3119: Pixel = 189;
			3120: Pixel = 190;
			3121: Pixel = 182;
			3122: Pixel = 176;
			3123: Pixel = 185;
			3124: Pixel = 184;
			3125: Pixel = 177;
			3126: Pixel = 171;
			3127: Pixel = 187;
			3128: Pixel = 193;
			3129: Pixel = 195;
			3130: Pixel = 195;
			3131: Pixel = 202;
			3132: Pixel = 205;
			3133: Pixel = 201;
			3134: Pixel = 200;
			3135: Pixel = 198;
			3136: Pixel = 201;
			3137: Pixel = 205;
			3138: Pixel = 199;
			3139: Pixel = 193;
			3140: Pixel = 207;
			3141: Pixel = 227;
			3142: Pixel = 176;
			3143: Pixel = 34;
			3144: Pixel = 46;
			3145: Pixel = 51;
			3146: Pixel = 48;
			3147: Pixel = 46;
			3148: Pixel = 53;
			3149: Pixel = 52;
			3150: Pixel = 106;
			3151: Pixel = 153;
			3152: Pixel = 145;
			3153: Pixel = 155;
			3154: Pixel = 161;
			3155: Pixel = 159;
			3156: Pixel = 158;
			3157: Pixel = 157;
			3158: Pixel = 157;
			3159: Pixel = 156;
			3160: Pixel = 155;
			3161: Pixel = 156;
			3162: Pixel = 97;
			3163: Pixel = 98;
			3164: Pixel = 97;
			3165: Pixel = 97;
			3166: Pixel = 97;
			3167: Pixel = 116;
			3168: Pixel = 147;
			3169: Pixel = 166;
			3170: Pixel = 172;
			3171: Pixel = 173;
			3172: Pixel = 170;
			3173: Pixel = 147;
			3174: Pixel = 106;
			3175: Pixel = 76;
			3176: Pixel = 87;
			3177: Pixel = 95;
			3178: Pixel = 98;
			3179: Pixel = 99;
			3180: Pixel = 98;
			3181: Pixel = 98;
			3182: Pixel = 99;
			3183: Pixel = 105;
			3184: Pixel = 96;
			3185: Pixel = 119;
			3186: Pixel = 205;
			3187: Pixel = 164;
			3188: Pixel = 140;
			3189: Pixel = 129;
			3190: Pixel = 111;
			3191: Pixel = 105;
			3192: Pixel = 106;
			3193: Pixel = 115;
			3194: Pixel = 113;
			3195: Pixel = 116;
			3196: Pixel = 140;
			3197: Pixel = 145;
			3198: Pixel = 141;
			3199: Pixel = 130;
			3200: Pixel = 140;
			3201: Pixel = 154;
			3202: Pixel = 149;
			3203: Pixel = 140;
			3204: Pixel = 153;
			3205: Pixel = 170;
			3206: Pixel = 160;
			3207: Pixel = 159;
			3208: Pixel = 177;
			3209: Pixel = 166;
			3210: Pixel = 169;
			3211: Pixel = 177;
			3212: Pixel = 172;
			3213: Pixel = 169;
			3214: Pixel = 169;
			3215: Pixel = 169;
			3216: Pixel = 176;
			3217: Pixel = 176;
			3218: Pixel = 181;
			3219: Pixel = 180;
			3220: Pixel = 186;
			3221: Pixel = 186;
			3222: Pixel = 178;
			3223: Pixel = 181;
			3224: Pixel = 175;
			3225: Pixel = 178;
			3226: Pixel = 170;
			3227: Pixel = 167;
			3228: Pixel = 185;
			3229: Pixel = 189;
			3230: Pixel = 186;
			3231: Pixel = 199;
			3232: Pixel = 204;
			3233: Pixel = 204;
			3234: Pixel = 196;
			3235: Pixel = 199;
			3236: Pixel = 199;
			3237: Pixel = 200;
			3238: Pixel = 203;
			3239: Pixel = 205;
			3240: Pixel = 169;
			3241: Pixel = 178;
			3242: Pixel = 196;
			3243: Pixel = 221;
			3244: Pixel = 122;
			3245: Pixel = 31;
			3246: Pixel = 49;
			3247: Pixel = 52;
			3248: Pixel = 48;
			3249: Pixel = 48;
			3250: Pixel = 49;
			3251: Pixel = 60;
			3252: Pixel = 141;
			3253: Pixel = 149;
			3254: Pixel = 150;
			3255: Pixel = 161;
			3256: Pixel = 160;
			3257: Pixel = 159;
			3258: Pixel = 159;
			3259: Pixel = 157;
			3260: Pixel = 158;
			3261: Pixel = 157;
			3262: Pixel = 157;
			3263: Pixel = 157;
			3264: Pixel = 97;
			3265: Pixel = 96;
			3266: Pixel = 96;
			3267: Pixel = 96;
			3268: Pixel = 97;
			3269: Pixel = 118;
			3270: Pixel = 151;
			3271: Pixel = 167;
			3272: Pixel = 171;
			3273: Pixel = 171;
			3274: Pixel = 168;
			3275: Pixel = 148;
			3276: Pixel = 105;
			3277: Pixel = 77;
			3278: Pixel = 87;
			3279: Pixel = 96;
			3280: Pixel = 99;
			3281: Pixel = 99;
			3282: Pixel = 98;
			3283: Pixel = 98;
			3284: Pixel = 99;
			3285: Pixel = 103;
			3286: Pixel = 94;
			3287: Pixel = 120;
			3288: Pixel = 201;
			3289: Pixel = 166;
			3290: Pixel = 151;
			3291: Pixel = 138;
			3292: Pixel = 122;
			3293: Pixel = 97;
			3294: Pixel = 103;
			3295: Pixel = 113;
			3296: Pixel = 112;
			3297: Pixel = 138;
			3298: Pixel = 139;
			3299: Pixel = 140;
			3300: Pixel = 125;
			3301: Pixel = 133;
			3302: Pixel = 152;
			3303: Pixel = 145;
			3304: Pixel = 146;
			3305: Pixel = 151;
			3306: Pixel = 149;
			3307: Pixel = 148;
			3308: Pixel = 158;
			3309: Pixel = 172;
			3310: Pixel = 166;
			3311: Pixel = 168;
			3312: Pixel = 166;
			3313: Pixel = 164;
			3314: Pixel = 167;
			3315: Pixel = 164;
			3316: Pixel = 164;
			3317: Pixel = 162;
			3318: Pixel = 164;
			3319: Pixel = 172;
			3320: Pixel = 174;
			3321: Pixel = 182;
			3322: Pixel = 179;
			3323: Pixel = 174;
			3324: Pixel = 171;
			3325: Pixel = 179;
			3326: Pixel = 171;
			3327: Pixel = 159;
			3328: Pixel = 177;
			3329: Pixel = 186;
			3330: Pixel = 190;
			3331: Pixel = 197;
			3332: Pixel = 203;
			3333: Pixel = 199;
			3334: Pixel = 193;
			3335: Pixel = 192;
			3336: Pixel = 198;
			3337: Pixel = 200;
			3338: Pixel = 200;
			3339: Pixel = 202;
			3340: Pixel = 209;
			3341: Pixel = 181;
			3342: Pixel = 160;
			3343: Pixel = 160;
			3344: Pixel = 163;
			3345: Pixel = 200;
			3346: Pixel = 63;
			3347: Pixel = 43;
			3348: Pixel = 55;
			3349: Pixel = 47;
			3350: Pixel = 46;
			3351: Pixel = 46;
			3352: Pixel = 59;
			3353: Pixel = 113;
			3354: Pixel = 152;
			3355: Pixel = 146;
			3356: Pixel = 157;
			3357: Pixel = 161;
			3358: Pixel = 159;
			3359: Pixel = 159;
			3360: Pixel = 158;
			3361: Pixel = 157;
			3362: Pixel = 156;
			3363: Pixel = 158;
			3364: Pixel = 157;
			3365: Pixel = 156;
			3366: Pixel = 97;
			3367: Pixel = 94;
			3368: Pixel = 94;
			3369: Pixel = 94;
			3370: Pixel = 96;
			3371: Pixel = 119;
			3372: Pixel = 151;
			3373: Pixel = 166;
			3374: Pixel = 170;
			3375: Pixel = 171;
			3376: Pixel = 168;
			3377: Pixel = 149;
			3378: Pixel = 106;
			3379: Pixel = 77;
			3380: Pixel = 87;
			3381: Pixel = 96;
			3382: Pixel = 99;
			3383: Pixel = 98;
			3384: Pixel = 97;
			3385: Pixel = 98;
			3386: Pixel = 100;
			3387: Pixel = 102;
			3388: Pixel = 87;
			3389: Pixel = 125;
			3390: Pixel = 198;
			3391: Pixel = 166;
			3392: Pixel = 151;
			3393: Pixel = 140;
			3394: Pixel = 126;
			3395: Pixel = 105;
			3396: Pixel = 103;
			3397: Pixel = 110;
			3398: Pixel = 141;
			3399: Pixel = 136;
			3400: Pixel = 133;
			3401: Pixel = 123;
			3402: Pixel = 132;
			3403: Pixel = 146;
			3404: Pixel = 143;
			3405: Pixel = 139;
			3406: Pixel = 140;
			3407: Pixel = 150;
			3408: Pixel = 146;
			3409: Pixel = 153;
			3410: Pixel = 162;
			3411: Pixel = 156;
			3412: Pixel = 164;
			3413: Pixel = 162;
			3414: Pixel = 164;
			3415: Pixel = 168;
			3416: Pixel = 162;
			3417: Pixel = 155;
			3418: Pixel = 161;
			3419: Pixel = 164;
			3420: Pixel = 165;
			3421: Pixel = 171;
			3422: Pixel = 167;
			3423: Pixel = 167;
			3424: Pixel = 170;
			3425: Pixel = 169;
			3426: Pixel = 166;
			3427: Pixel = 158;
			3428: Pixel = 169;
			3429: Pixel = 180;
			3430: Pixel = 183;
			3431: Pixel = 190;
			3432: Pixel = 200;
			3433: Pixel = 201;
			3434: Pixel = 193;
			3435: Pixel = 192;
			3436: Pixel = 192;
			3437: Pixel = 197;
			3438: Pixel = 201;
			3439: Pixel = 201;
			3440: Pixel = 201;
			3441: Pixel = 208;
			3442: Pixel = 201;
			3443: Pixel = 160;
			3444: Pixel = 168;
			3445: Pixel = 149;
			3446: Pixel = 179;
			3447: Pixel = 166;
			3448: Pixel = 34;
			3449: Pixel = 46;
			3450: Pixel = 52;
			3451: Pixel = 44;
			3452: Pixel = 49;
			3453: Pixel = 48;
			3454: Pixel = 83;
			3455: Pixel = 148;
			3456: Pixel = 147;
			3457: Pixel = 150;
			3458: Pixel = 161;
			3459: Pixel = 160;
			3460: Pixel = 157;
			3461: Pixel = 157;
			3462: Pixel = 158;
			3463: Pixel = 157;
			3464: Pixel = 156;
			3465: Pixel = 157;
			3466: Pixel = 156;
			3467: Pixel = 156;
			3468: Pixel = 96;
			3469: Pixel = 96;
			3470: Pixel = 95;
			3471: Pixel = 95;
			3472: Pixel = 100;
			3473: Pixel = 122;
			3474: Pixel = 150;
			3475: Pixel = 167;
			3476: Pixel = 171;
			3477: Pixel = 172;
			3478: Pixel = 169;
			3479: Pixel = 151;
			3480: Pixel = 109;
			3481: Pixel = 76;
			3482: Pixel = 86;
			3483: Pixel = 95;
			3484: Pixel = 97;
			3485: Pixel = 96;
			3486: Pixel = 97;
			3487: Pixel = 97;
			3488: Pixel = 98;
			3489: Pixel = 101;
			3490: Pixel = 83;
			3491: Pixel = 134;
			3492: Pixel = 206;
			3493: Pixel = 176;
			3494: Pixel = 159;
			3495: Pixel = 145;
			3496: Pixel = 138;
			3497: Pixel = 110;
			3498: Pixel = 104;
			3499: Pixel = 135;
			3500: Pixel = 134;
			3501: Pixel = 135;
			3502: Pixel = 120;
			3503: Pixel = 129;
			3504: Pixel = 145;
			3505: Pixel = 144;
			3506: Pixel = 133;
			3507: Pixel = 131;
			3508: Pixel = 149;
			3509: Pixel = 139;
			3510: Pixel = 153;
			3511: Pixel = 161;
			3512: Pixel = 146;
			3513: Pixel = 153;
			3514: Pixel = 157;
			3515: Pixel = 144;
			3516: Pixel = 138;
			3517: Pixel = 138;
			3518: Pixel = 159;
			3519: Pixel = 162;
			3520: Pixel = 163;
			3521: Pixel = 161;
			3522: Pixel = 165;
			3523: Pixel = 163;
			3524: Pixel = 166;
			3525: Pixel = 166;
			3526: Pixel = 161;
			3527: Pixel = 156;
			3528: Pixel = 157;
			3529: Pixel = 173;
			3530: Pixel = 181;
			3531: Pixel = 184;
			3532: Pixel = 196;
			3533: Pixel = 195;
			3534: Pixel = 188;
			3535: Pixel = 187;
			3536: Pixel = 192;
			3537: Pixel = 196;
			3538: Pixel = 198;
			3539: Pixel = 202;
			3540: Pixel = 203;
			3541: Pixel = 202;
			3542: Pixel = 203;
			3543: Pixel = 212;
			3544: Pixel = 177;
			3545: Pixel = 161;
			3546: Pixel = 148;
			3547: Pixel = 129;
			3548: Pixel = 196;
			3549: Pixel = 115;
			3550: Pixel = 30;
			3551: Pixel = 54;
			3552: Pixel = 49;
			3553: Pixel = 55;
			3554: Pixel = 53;
			3555: Pixel = 53;
			3556: Pixel = 118;
			3557: Pixel = 154;
			3558: Pixel = 145;
			3559: Pixel = 157;
			3560: Pixel = 159;
			3561: Pixel = 157;
			3562: Pixel = 156;
			3563: Pixel = 156;
			3564: Pixel = 157;
			3565: Pixel = 156;
			3566: Pixel = 156;
			3567: Pixel = 157;
			3568: Pixel = 156;
			3569: Pixel = 156;
			3570: Pixel = 97;
			3571: Pixel = 98;
			3572: Pixel = 97;
			3573: Pixel = 99;
			3574: Pixel = 104;
			3575: Pixel = 122;
			3576: Pixel = 150;
			3577: Pixel = 167;
			3578: Pixel = 172;
			3579: Pixel = 172;
			3580: Pixel = 170;
			3581: Pixel = 152;
			3582: Pixel = 107;
			3583: Pixel = 73;
			3584: Pixel = 83;
			3585: Pixel = 95;
			3586: Pixel = 98;
			3587: Pixel = 96;
			3588: Pixel = 97;
			3589: Pixel = 98;
			3590: Pixel = 98;
			3591: Pixel = 100;
			3592: Pixel = 80;
			3593: Pixel = 135;
			3594: Pixel = 213;
			3595: Pixel = 181;
			3596: Pixel = 164;
			3597: Pixel = 154;
			3598: Pixel = 151;
			3599: Pixel = 118;
			3600: Pixel = 118;
			3601: Pixel = 130;
			3602: Pixel = 132;
			3603: Pixel = 119;
			3604: Pixel = 128;
			3605: Pixel = 143;
			3606: Pixel = 138;
			3607: Pixel = 130;
			3608: Pixel = 128;
			3609: Pixel = 142;
			3610: Pixel = 137;
			3611: Pixel = 146;
			3612: Pixel = 148;
			3613: Pixel = 124;
			3614: Pixel = 127;
			3615: Pixel = 113;
			3616: Pixel = 116;
			3617: Pixel = 124;
			3618: Pixel = 151;
			3619: Pixel = 120;
			3620: Pixel = 137;
			3621: Pixel = 152;
			3622: Pixel = 153;
			3623: Pixel = 155;
			3624: Pixel = 152;
			3625: Pixel = 157;
			3626: Pixel = 134;
			3627: Pixel = 126;
			3628: Pixel = 151;
			3629: Pixel = 155;
			3630: Pixel = 177;
			3631: Pixel = 179;
			3632: Pixel = 191;
			3633: Pixel = 199;
			3634: Pixel = 195;
			3635: Pixel = 189;
			3636: Pixel = 190;
			3637: Pixel = 194;
			3638: Pixel = 198;
			3639: Pixel = 199;
			3640: Pixel = 201;
			3641: Pixel = 203;
			3642: Pixel = 201;
			3643: Pixel = 202;
			3644: Pixel = 215;
			3645: Pixel = 204;
			3646: Pixel = 154;
			3647: Pixel = 115;
			3648: Pixel = 87;
			3649: Pixel = 141;
			3650: Pixel = 209;
			3651: Pixel = 53;
			3652: Pixel = 37;
			3653: Pixel = 51;
			3654: Pixel = 46;
			3655: Pixel = 55;
			3656: Pixel = 51;
			3657: Pixel = 74;
			3658: Pixel = 146;
			3659: Pixel = 148;
			3660: Pixel = 152;
			3661: Pixel = 159;
			3662: Pixel = 159;
			3663: Pixel = 157;
			3664: Pixel = 156;
			3665: Pixel = 155;
			3666: Pixel = 156;
			3667: Pixel = 155;
			3668: Pixel = 155;
			3669: Pixel = 156;
			3670: Pixel = 154;
			3671: Pixel = 153;
			3672: Pixel = 99;
			3673: Pixel = 98;
			3674: Pixel = 98;
			3675: Pixel = 100;
			3676: Pixel = 105;
			3677: Pixel = 126;
			3678: Pixel = 151;
			3679: Pixel = 168;
			3680: Pixel = 173;
			3681: Pixel = 173;
			3682: Pixel = 171;
			3683: Pixel = 152;
			3684: Pixel = 107;
			3685: Pixel = 72;
			3686: Pixel = 82;
			3687: Pixel = 94;
			3688: Pixel = 97;
			3689: Pixel = 99;
			3690: Pixel = 99;
			3691: Pixel = 99;
			3692: Pixel = 99;
			3693: Pixel = 100;
			3694: Pixel = 80;
			3695: Pixel = 131;
			3696: Pixel = 212;
			3697: Pixel = 189;
			3698: Pixel = 171;
			3699: Pixel = 143;
			3700: Pixel = 150;
			3701: Pixel = 125;
			3702: Pixel = 115;
			3703: Pixel = 124;
			3704: Pixel = 116;
			3705: Pixel = 122;
			3706: Pixel = 140;
			3707: Pixel = 137;
			3708: Pixel = 126;
			3709: Pixel = 125;
			3710: Pixel = 135;
			3711: Pixel = 133;
			3712: Pixel = 139;
			3713: Pixel = 147;
			3714: Pixel = 127;
			3715: Pixel = 131;
			3716: Pixel = 118;
			3717: Pixel = 103;
			3718: Pixel = 77;
			3719: Pixel = 96;
			3720: Pixel = 168;
			3721: Pixel = 146;
			3722: Pixel = 111;
			3723: Pixel = 96;
			3724: Pixel = 101;
			3725: Pixel = 105;
			3726: Pixel = 88;
			3727: Pixel = 73;
			3728: Pixel = 65;
			3729: Pixel = 46;
			3730: Pixel = 150;
			3731: Pixel = 173;
			3732: Pixel = 172;
			3733: Pixel = 192;
			3734: Pixel = 199;
			3735: Pixel = 193;
			3736: Pixel = 195;
			3737: Pixel = 193;
			3738: Pixel = 192;
			3739: Pixel = 197;
			3740: Pixel = 200;
			3741: Pixel = 200;
			3742: Pixel = 200;
			3743: Pixel = 204;
			3744: Pixel = 210;
			3745: Pixel = 209;
			3746: Pixel = 186;
			3747: Pixel = 135;
			3748: Pixel = 91;
			3749: Pixel = 79;
			3750: Pixel = 118;
			3751: Pixel = 219;
			3752: Pixel = 129;
			3753: Pixel = 28;
			3754: Pixel = 51;
			3755: Pixel = 46;
			3756: Pixel = 45;
			3757: Pixel = 52;
			3758: Pixel = 47;
			3759: Pixel = 113;
			3760: Pixel = 152;
			3761: Pixel = 145;
			3762: Pixel = 159;
			3763: Pixel = 160;
			3764: Pixel = 159;
			3765: Pixel = 158;
			3766: Pixel = 156;
			3767: Pixel = 156;
			3768: Pixel = 155;
			3769: Pixel = 154;
			3770: Pixel = 154;
			3771: Pixel = 153;
			3772: Pixel = 154;
			3773: Pixel = 153;
			3774: Pixel = 99;
			3775: Pixel = 102;
			3776: Pixel = 98;
			3777: Pixel = 101;
			3778: Pixel = 108;
			3779: Pixel = 126;
			3780: Pixel = 153;
			3781: Pixel = 169;
			3782: Pixel = 172;
			3783: Pixel = 173;
			3784: Pixel = 171;
			3785: Pixel = 153;
			3786: Pixel = 108;
			3787: Pixel = 73;
			3788: Pixel = 83;
			3789: Pixel = 94;
			3790: Pixel = 97;
			3791: Pixel = 98;
			3792: Pixel = 99;
			3793: Pixel = 99;
			3794: Pixel = 99;
			3795: Pixel = 101;
			3796: Pixel = 86;
			3797: Pixel = 113;
			3798: Pixel = 209;
			3799: Pixel = 199;
			3800: Pixel = 180;
			3801: Pixel = 126;
			3802: Pixel = 130;
			3803: Pixel = 117;
			3804: Pixel = 116;
			3805: Pixel = 114;
			3806: Pixel = 114;
			3807: Pixel = 138;
			3808: Pixel = 135;
			3809: Pixel = 125;
			3810: Pixel = 127;
			3811: Pixel = 135;
			3812: Pixel = 128;
			3813: Pixel = 134;
			3814: Pixel = 143;
			3815: Pixel = 118;
			3816: Pixel = 131;
			3817: Pixel = 125;
			3818: Pixel = 112;
			3819: Pixel = 111;
			3820: Pixel = 97;
			3821: Pixel = 83;
			3822: Pixel = 109;
			3823: Pixel = 111;
			3824: Pixel = 76;
			3825: Pixel = 81;
			3826: Pixel = 81;
			3827: Pixel = 66;
			3828: Pixel = 53;
			3829: Pixel = 30;
			3830: Pixel = 42;
			3831: Pixel = 124;
			3832: Pixel = 158;
			3833: Pixel = 179;
			3834: Pixel = 202;
			3835: Pixel = 197;
			3836: Pixel = 192;
			3837: Pixel = 193;
			3838: Pixel = 195;
			3839: Pixel = 191;
			3840: Pixel = 193;
			3841: Pixel = 197;
			3842: Pixel = 198;
			3843: Pixel = 197;
			3844: Pixel = 208;
			3845: Pixel = 207;
			3846: Pixel = 169;
			3847: Pixel = 120;
			3848: Pixel = 89;
			3849: Pixel = 83;
			3850: Pixel = 91;
			3851: Pixel = 129;
			3852: Pixel = 194;
			3853: Pixel = 159;
			3854: Pixel = 45;
			3855: Pixel = 45;
			3856: Pixel = 51;
			3857: Pixel = 48;
			3858: Pixel = 52;
			3859: Pixel = 44;
			3860: Pixel = 59;
			3861: Pixel = 143;
			3862: Pixel = 145;
			3863: Pixel = 153;
			3864: Pixel = 163;
			3865: Pixel = 159;
			3866: Pixel = 160;
			3867: Pixel = 159;
			3868: Pixel = 157;
			3869: Pixel = 156;
			3870: Pixel = 154;
			3871: Pixel = 154;
			3872: Pixel = 154;
			3873: Pixel = 154;
			3874: Pixel = 153;
			3875: Pixel = 153;
			3876: Pixel = 103;
			3877: Pixel = 103;
			3878: Pixel = 97;
			3879: Pixel = 99;
			3880: Pixel = 108;
			3881: Pixel = 126;
			3882: Pixel = 151;
			3883: Pixel = 169;
			3884: Pixel = 171;
			3885: Pixel = 172;
			3886: Pixel = 170;
			3887: Pixel = 153;
			3888: Pixel = 107;
			3889: Pixel = 74;
			3890: Pixel = 84;
			3891: Pixel = 95;
			3892: Pixel = 97;
			3893: Pixel = 97;
			3894: Pixel = 100;
			3895: Pixel = 99;
			3896: Pixel = 99;
			3897: Pixel = 97;
			3898: Pixel = 91;
			3899: Pixel = 93;
			3900: Pixel = 199;
			3901: Pixel = 205;
			3902: Pixel = 181;
			3903: Pixel = 126;
			3904: Pixel = 140;
			3905: Pixel = 138;
			3906: Pixel = 112;
			3907: Pixel = 109;
			3908: Pixel = 134;
			3909: Pixel = 138;
			3910: Pixel = 124;
			3911: Pixel = 122;
			3912: Pixel = 134;
			3913: Pixel = 129;
			3914: Pixel = 131;
			3915: Pixel = 138;
			3916: Pixel = 118;
			3917: Pixel = 131;
			3918: Pixel = 127;
			3919: Pixel = 101;
			3920: Pixel = 102;
			3921: Pixel = 76;
			3922: Pixel = 56;
			3923: Pixel = 63;
			3924: Pixel = 106;
			3925: Pixel = 94;
			3926: Pixel = 88;
			3927: Pixel = 105;
			3928: Pixel = 71;
			3929: Pixel = 75;
			3930: Pixel = 42;
			3931: Pixel = 46;
			3932: Pixel = 135;
			3933: Pixel = 150;
			3934: Pixel = 178;
			3935: Pixel = 190;
			3936: Pixel = 190;
			3937: Pixel = 193;
			3938: Pixel = 190;
			3939: Pixel = 189;
			3940: Pixel = 192;
			3941: Pixel = 191;
			3942: Pixel = 192;
			3943: Pixel = 193;
			3944: Pixel = 202;
			3945: Pixel = 206;
			3946: Pixel = 187;
			3947: Pixel = 135;
			3948: Pixel = 80;
			3949: Pixel = 80;
			3950: Pixel = 95;
			3951: Pixel = 125;
			3952: Pixel = 148;
			3953: Pixel = 205;
			3954: Pixel = 144;
			3955: Pixel = 32;
			3956: Pixel = 44;
			3957: Pixel = 53;
			3958: Pixel = 45;
			3959: Pixel = 46;
			3960: Pixel = 58;
			3961: Pixel = 46;
			3962: Pixel = 96;
			3963: Pixel = 152;
			3964: Pixel = 146;
			3965: Pixel = 162;
			3966: Pixel = 163;
			3967: Pixel = 160;
			3968: Pixel = 160;
			3969: Pixel = 159;
			3970: Pixel = 158;
			3971: Pixel = 157;
			3972: Pixel = 156;
			3973: Pixel = 155;
			3974: Pixel = 154;
			3975: Pixel = 154;
			3976: Pixel = 154;
			3977: Pixel = 152;
			3978: Pixel = 106;
			3979: Pixel = 103;
			3980: Pixel = 101;
			3981: Pixel = 100;
			3982: Pixel = 104;
			3983: Pixel = 125;
			3984: Pixel = 151;
			3985: Pixel = 167;
			3986: Pixel = 170;
			3987: Pixel = 170;
			3988: Pixel = 169;
			3989: Pixel = 153;
			3990: Pixel = 109;
			3991: Pixel = 74;
			3992: Pixel = 83;
			3993: Pixel = 93;
			3994: Pixel = 96;
			3995: Pixel = 98;
			3996: Pixel = 99;
			3997: Pixel = 98;
			3998: Pixel = 98;
			3999: Pixel = 98;
			4000: Pixel = 100;
			4001: Pixel = 79;
			4002: Pixel = 171;
			4003: Pixel = 205;
			4004: Pixel = 186;
			4005: Pixel = 145;
			4006: Pixel = 141;
			4007: Pixel = 137;
			4008: Pixel = 106;
			4009: Pixel = 129;
			4010: Pixel = 136;
			4011: Pixel = 121;
			4012: Pixel = 122;
			4013: Pixel = 130;
			4014: Pixel = 127;
			4015: Pixel = 124;
			4016: Pixel = 139;
			4017: Pixel = 138;
			4018: Pixel = 119;
			4019: Pixel = 119;
			4020: Pixel = 76;
			4021: Pixel = 77;
			4022: Pixel = 68;
			4023: Pixel = 55;
			4024: Pixel = 46;
			4025: Pixel = 105;
			4026: Pixel = 101;
			4027: Pixel = 49;
			4028: Pixel = 83;
			4029: Pixel = 88;
			4030: Pixel = 56;
			4031: Pixel = 62;
			4032: Pixel = 66;
			4033: Pixel = 136;
			4034: Pixel = 152;
			4035: Pixel = 179;
			4036: Pixel = 189;
			4037: Pixel = 178;
			4038: Pixel = 186;
			4039: Pixel = 187;
			4040: Pixel = 186;
			4041: Pixel = 186;
			4042: Pixel = 190;
			4043: Pixel = 190;
			4044: Pixel = 194;
			4045: Pixel = 207;
			4046: Pixel = 185;
			4047: Pixel = 127;
			4048: Pixel = 103;
			4049: Pixel = 130;
			4050: Pixel = 124;
			4051: Pixel = 137;
			4052: Pixel = 158;
			4053: Pixel = 163;
			4054: Pixel = 196;
			4055: Pixel = 150;
			4056: Pixel = 38;
			4057: Pixel = 48;
			4058: Pixel = 55;
			4059: Pixel = 52;
			4060: Pixel = 45;
			4061: Pixel = 49;
			4062: Pixel = 55;
			4063: Pixel = 58;
			4064: Pixel = 134;
			4065: Pixel = 147;
			4066: Pixel = 153;
			4067: Pixel = 165;
			4068: Pixel = 163;
			4069: Pixel = 162;
			4070: Pixel = 161;
			4071: Pixel = 160;
			4072: Pixel = 158;
			4073: Pixel = 158;
			4074: Pixel = 155;
			4075: Pixel = 155;
			4076: Pixel = 155;
			4077: Pixel = 155;
			4078: Pixel = 154;
			4079: Pixel = 151;
			4080: Pixel = 106;
			4081: Pixel = 104;
			4082: Pixel = 102;
			4083: Pixel = 100;
			4084: Pixel = 103;
			4085: Pixel = 123;
			4086: Pixel = 150;
			4087: Pixel = 168;
			4088: Pixel = 171;
			4089: Pixel = 171;
			4090: Pixel = 170;
			4091: Pixel = 153;
			4092: Pixel = 111;
			4093: Pixel = 73;
			4094: Pixel = 84;
			4095: Pixel = 93;
			4096: Pixel = 95;
			4097: Pixel = 97;
			4098: Pixel = 99;
			4099: Pixel = 98;
			4100: Pixel = 97;
			4101: Pixel = 98;
			4102: Pixel = 104;
			4103: Pixel = 82;
			4104: Pixel = 137;
			4105: Pixel = 213;
			4106: Pixel = 191;
			4107: Pixel = 170;
			4108: Pixel = 153;
			4109: Pixel = 113;
			4110: Pixel = 120;
			4111: Pixel = 139;
			4112: Pixel = 122;
			4113: Pixel = 114;
			4114: Pixel = 127;
			4115: Pixel = 124;
			4116: Pixel = 122;
			4117: Pixel = 133;
			4118: Pixel = 111;
			4119: Pixel = 124;
			4120: Pixel = 105;
			4121: Pixel = 68;
			4122: Pixel = 75;
			4123: Pixel = 63;
			4124: Pixel = 54;
			4125: Pixel = 43;
			4126: Pixel = 67;
			4127: Pixel = 94;
			4128: Pixel = 51;
			4129: Pixel = 87;
			4130: Pixel = 106;
			4131: Pixel = 66;
			4132: Pixel = 45;
			4133: Pixel = 94;
			4134: Pixel = 143;
			4135: Pixel = 147;
			4136: Pixel = 186;
			4137: Pixel = 193;
			4138: Pixel = 177;
			4139: Pixel = 182;
			4140: Pixel = 182;
			4141: Pixel = 178;
			4142: Pixel = 179;
			4143: Pixel = 187;
			4144: Pixel = 190;
			4145: Pixel = 192;
			4146: Pixel = 195;
			4147: Pixel = 138;
			4148: Pixel = 78;
			4149: Pixel = 98;
			4150: Pixel = 110;
			4151: Pixel = 139;
			4152: Pixel = 168;
			4153: Pixel = 170;
			4154: Pixel = 168;
			4155: Pixel = 196;
			4156: Pixel = 160;
			4157: Pixel = 41;
			4158: Pixel = 41;
			4159: Pixel = 53;
			4160: Pixel = 54;
			4161: Pixel = 51;
			4162: Pixel = 46;
			4163: Pixel = 53;
			4164: Pixel = 44;
			4165: Pixel = 84;
			4166: Pixel = 149;
			4167: Pixel = 144;
			4168: Pixel = 162;
			4169: Pixel = 165;
			4170: Pixel = 164;
			4171: Pixel = 164;
			4172: Pixel = 162;
			4173: Pixel = 161;
			4174: Pixel = 158;
			4175: Pixel = 158;
			4176: Pixel = 156;
			4177: Pixel = 156;
			4178: Pixel = 155;
			4179: Pixel = 154;
			4180: Pixel = 153;
			4181: Pixel = 152;
			4182: Pixel = 107;
			4183: Pixel = 106;
			4184: Pixel = 102;
			4185: Pixel = 99;
			4186: Pixel = 100;
			4187: Pixel = 120;
			4188: Pixel = 150;
			4189: Pixel = 169;
			4190: Pixel = 171;
			4191: Pixel = 172;
			4192: Pixel = 170;
			4193: Pixel = 154;
			4194: Pixel = 112;
			4195: Pixel = 71;
			4196: Pixel = 83;
			4197: Pixel = 92;
			4198: Pixel = 95;
			4199: Pixel = 96;
			4200: Pixel = 97;
			4201: Pixel = 96;
			4202: Pixel = 97;
			4203: Pixel = 101;
			4204: Pixel = 106;
			4205: Pixel = 99;
			4206: Pixel = 94;
			4207: Pixel = 199;
			4208: Pixel = 199;
			4209: Pixel = 171;
			4210: Pixel = 160;
			4211: Pixel = 111;
			4212: Pixel = 134;
			4213: Pixel = 123;
			4214: Pixel = 115;
			4215: Pixel = 130;
			4216: Pixel = 122;
			4217: Pixel = 121;
			4218: Pixel = 131;
			4219: Pixel = 132;
			4220: Pixel = 101;
			4221: Pixel = 72;
			4222: Pixel = 72;
			4223: Pixel = 79;
			4224: Pixel = 62;
			4225: Pixel = 61;
			4226: Pixel = 76;
			4227: Pixel = 37;
			4228: Pixel = 84;
			4229: Pixel = 51;
			4230: Pixel = 55;
			4231: Pixel = 76;
			4232: Pixel = 72;
			4233: Pixel = 83;
			4234: Pixel = 79;
			4235: Pixel = 125;
			4236: Pixel = 145;
			4237: Pixel = 191;
			4238: Pixel = 196;
			4239: Pixel = 184;
			4240: Pixel = 180;
			4241: Pixel = 182;
			4242: Pixel = 176;
			4243: Pixel = 174;
			4244: Pixel = 178;
			4245: Pixel = 188;
			4246: Pixel = 189;
			4247: Pixel = 192;
			4248: Pixel = 151;
			4249: Pixel = 61;
			4250: Pixel = 87;
			4251: Pixel = 108;
			4252: Pixel = 124;
			4253: Pixel = 120;
			4254: Pixel = 154;
			4255: Pixel = 172;
			4256: Pixel = 196;
			4257: Pixel = 135;
			4258: Pixel = 41;
			4259: Pixel = 40;
			4260: Pixel = 51;
			4261: Pixel = 53;
			4262: Pixel = 56;
			4263: Pixel = 50;
			4264: Pixel = 46;
			4265: Pixel = 51;
			4266: Pixel = 53;
			4267: Pixel = 114;
			4268: Pixel = 140;
			4269: Pixel = 148;
			4270: Pixel = 167;
			4271: Pixel = 165;
			4272: Pixel = 164;
			4273: Pixel = 163;
			4274: Pixel = 163;
			4275: Pixel = 162;
			4276: Pixel = 160;
			4277: Pixel = 158;
			4278: Pixel = 157;
			4279: Pixel = 157;
			4280: Pixel = 156;
			4281: Pixel = 155;
			4282: Pixel = 153;
			4283: Pixel = 151;
			4284: Pixel = 108;
			4285: Pixel = 106;
			4286: Pixel = 103;
			4287: Pixel = 99;
			4288: Pixel = 95;
			4289: Pixel = 116;
			4290: Pixel = 149;
			4291: Pixel = 168;
			4292: Pixel = 172;
			4293: Pixel = 173;
			4294: Pixel = 171;
			4295: Pixel = 154;
			4296: Pixel = 110;
			4297: Pixel = 72;
			4298: Pixel = 81;
			4299: Pixel = 90;
			4300: Pixel = 96;
			4301: Pixel = 97;
			4302: Pixel = 97;
			4303: Pixel = 98;
			4304: Pixel = 98;
			4305: Pixel = 102;
			4306: Pixel = 106;
			4307: Pixel = 109;
			4308: Pixel = 87;
			4309: Pixel = 131;
			4310: Pixel = 210;
			4311: Pixel = 189;
			4312: Pixel = 152;
			4313: Pixel = 125;
			4314: Pixel = 125;
			4315: Pixel = 118;
			4316: Pixel = 127;
			4317: Pixel = 128;
			4318: Pixel = 122;
			4319: Pixel = 125;
			4320: Pixel = 125;
			4321: Pixel = 109;
			4322: Pixel = 89;
			4323: Pixel = 81;
			4324: Pixel = 87;
			4325: Pixel = 70;
			4326: Pixel = 33;
			4327: Pixel = 82;
			4328: Pixel = 66;
			4329: Pixel = 51;
			4330: Pixel = 67;
			4331: Pixel = 57;
			4332: Pixel = 65;
			4333: Pixel = 67;
			4334: Pixel = 72;
			4335: Pixel = 102;
			4336: Pixel = 122;
			4337: Pixel = 124;
			4338: Pixel = 188;
			4339: Pixel = 194;
			4340: Pixel = 187;
			4341: Pixel = 180;
			4342: Pixel = 178;
			4343: Pixel = 179;
			4344: Pixel = 172;
			4345: Pixel = 178;
			4346: Pixel = 182;
			4347: Pixel = 184;
			4348: Pixel = 184;
			4349: Pixel = 194;
			4350: Pixel = 178;
			4351: Pixel = 102;
			4352: Pixel = 92;
			4353: Pixel = 102;
			4354: Pixel = 117;
			4355: Pixel = 125;
			4356: Pixel = 155;
			4357: Pixel = 181;
			4358: Pixel = 106;
			4359: Pixel = 35;
			4360: Pixel = 42;
			4361: Pixel = 52;
			4362: Pixel = 53;
			4363: Pixel = 54;
			4364: Pixel = 54;
			4365: Pixel = 45;
			4366: Pixel = 49;
			4367: Pixel = 51;
			4368: Pixel = 74;
			4369: Pixel = 129;
			4370: Pixel = 128;
			4371: Pixel = 159;
			4372: Pixel = 169;
			4373: Pixel = 163;
			4374: Pixel = 162;
			4375: Pixel = 162;
			4376: Pixel = 163;
			4377: Pixel = 162;
			4378: Pixel = 160;
			4379: Pixel = 159;
			4380: Pixel = 159;
			4381: Pixel = 158;
			4382: Pixel = 156;
			4383: Pixel = 155;
			4384: Pixel = 154;
			4385: Pixel = 151;
			4386: Pixel = 108;
			4387: Pixel = 105;
			4388: Pixel = 102;
			4389: Pixel = 100;
			4390: Pixel = 92;
			4391: Pixel = 112;
			4392: Pixel = 148;
			4393: Pixel = 167;
			4394: Pixel = 172;
			4395: Pixel = 173;
			4396: Pixel = 173;
			4397: Pixel = 155;
			4398: Pixel = 113;
			4399: Pixel = 70;
			4400: Pixel = 79;
			4401: Pixel = 89;
			4402: Pixel = 96;
			4403: Pixel = 97;
			4404: Pixel = 96;
			4405: Pixel = 97;
			4406: Pixel = 98;
			4407: Pixel = 103;
			4408: Pixel = 108;
			4409: Pixel = 112;
			4410: Pixel = 102;
			4411: Pixel = 96;
			4412: Pixel = 202;
			4413: Pixel = 205;
			4414: Pixel = 162;
			4415: Pixel = 122;
			4416: Pixel = 111;
			4417: Pixel = 118;
			4418: Pixel = 126;
			4419: Pixel = 115;
			4420: Pixel = 128;
			4421: Pixel = 122;
			4422: Pixel = 125;
			4423: Pixel = 85;
			4424: Pixel = 62;
			4425: Pixel = 70;
			4426: Pixel = 88;
			4427: Pixel = 63;
			4428: Pixel = 50;
			4429: Pixel = 72;
			4430: Pixel = 80;
			4431: Pixel = 56;
			4432: Pixel = 44;
			4433: Pixel = 53;
			4434: Pixel = 59;
			4435: Pixel = 54;
			4436: Pixel = 82;
			4437: Pixel = 86;
			4438: Pixel = 122;
			4439: Pixel = 163;
			4440: Pixel = 179;
			4441: Pixel = 181;
			4442: Pixel = 178;
			4443: Pixel = 171;
			4444: Pixel = 174;
			4445: Pixel = 175;
			4446: Pixel = 174;
			4447: Pixel = 173;
			4448: Pixel = 187;
			4449: Pixel = 193;
			4450: Pixel = 194;
			4451: Pixel = 198;
			4452: Pixel = 198;
			4453: Pixel = 140;
			4454: Pixel = 76;
			4455: Pixel = 82;
			4456: Pixel = 90;
			4457: Pixel = 129;
			4458: Pixel = 154;
			4459: Pixel = 111;
			4460: Pixel = 32;
			4461: Pixel = 44;
			4462: Pixel = 49;
			4463: Pixel = 54;
			4464: Pixel = 57;
			4465: Pixel = 57;
			4466: Pixel = 49;
			4467: Pixel = 44;
			4468: Pixel = 52;
			4469: Pixel = 51;
			4470: Pixel = 101;
			4471: Pixel = 131;
			4472: Pixel = 131;
			4473: Pixel = 166;
			4474: Pixel = 166;
			4475: Pixel = 164;
			4476: Pixel = 163;
			4477: Pixel = 163;
			4478: Pixel = 163;
			4479: Pixel = 161;
			4480: Pixel = 161;
			4481: Pixel = 160;
			4482: Pixel = 160;
			4483: Pixel = 157;
			4484: Pixel = 157;
			4485: Pixel = 156;
			4486: Pixel = 153;
			4487: Pixel = 152;
			4488: Pixel = 105;
			4489: Pixel = 105;
			4490: Pixel = 103;
			4491: Pixel = 98;
			4492: Pixel = 90;
			4493: Pixel = 110;
			4494: Pixel = 146;
			4495: Pixel = 166;
			4496: Pixel = 172;
			4497: Pixel = 173;
			4498: Pixel = 172;
			4499: Pixel = 155;
			4500: Pixel = 113;
			4501: Pixel = 71;
			4502: Pixel = 81;
			4503: Pixel = 92;
			4504: Pixel = 97;
			4505: Pixel = 99;
			4506: Pixel = 99;
			4507: Pixel = 97;
			4508: Pixel = 98;
			4509: Pixel = 103;
			4510: Pixel = 110;
			4511: Pixel = 113;
			4512: Pixel = 106;
			4513: Pixel = 98;
			4514: Pixel = 202;
			4515: Pixel = 214;
			4516: Pixel = 135;
			4517: Pixel = 115;
			4518: Pixel = 122;
			4519: Pixel = 116;
			4520: Pixel = 116;
			4521: Pixel = 136;
			4522: Pixel = 134;
			4523: Pixel = 102;
			4524: Pixel = 73;
			4525: Pixel = 75;
			4526: Pixel = 55;
			4527: Pixel = 45;
			4528: Pixel = 72;
			4529: Pixel = 77;
			4530: Pixel = 64;
			4531: Pixel = 54;
			4532: Pixel = 100;
			4533: Pixel = 71;
			4534: Pixel = 45;
			4535: Pixel = 48;
			4536: Pixel = 32;
			4537: Pixel = 65;
			4538: Pixel = 101;
			4539: Pixel = 112;
			4540: Pixel = 159;
			4541: Pixel = 179;
			4542: Pixel = 184;
			4543: Pixel = 183;
			4544: Pixel = 164;
			4545: Pixel = 167;
			4546: Pixel = 179;
			4547: Pixel = 166;
			4548: Pixel = 169;
			4549: Pixel = 184;
			4550: Pixel = 198;
			4551: Pixel = 199;
			4552: Pixel = 196;
			4553: Pixel = 198;
			4554: Pixel = 199;
			4555: Pixel = 159;
			4556: Pixel = 86;
			4557: Pixel = 50;
			4558: Pixel = 75;
			4559: Pixel = 112;
			4560: Pixel = 154;
			4561: Pixel = 98;
			4562: Pixel = 42;
			4563: Pixel = 44;
			4564: Pixel = 50;
			4565: Pixel = 56;
			4566: Pixel = 59;
			4567: Pixel = 58;
			4568: Pixel = 47;
			4569: Pixel = 45;
			4570: Pixel = 47;
			4571: Pixel = 60;
			4572: Pixel = 128;
			4573: Pixel = 129;
			4574: Pixel = 143;
			4575: Pixel = 162;
			4576: Pixel = 166;
			4577: Pixel = 165;
			4578: Pixel = 164;
			4579: Pixel = 161;
			4580: Pixel = 162;
			4581: Pixel = 162;
			4582: Pixel = 162;
			4583: Pixel = 160;
			4584: Pixel = 160;
			4585: Pixel = 158;
			4586: Pixel = 158;
			4587: Pixel = 157;
			4588: Pixel = 154;
			4589: Pixel = 151;
			4590: Pixel = 104;
			4591: Pixel = 105;
			4592: Pixel = 102;
			4593: Pixel = 99;
			4594: Pixel = 91;
			4595: Pixel = 110;
			4596: Pixel = 147;
			4597: Pixel = 166;
			4598: Pixel = 172;
			4599: Pixel = 173;
			4600: Pixel = 171;
			4601: Pixel = 156;
			4602: Pixel = 114;
			4603: Pixel = 73;
			4604: Pixel = 81;
			4605: Pixel = 93;
			4606: Pixel = 97;
			4607: Pixel = 99;
			4608: Pixel = 101;
			4609: Pixel = 99;
			4610: Pixel = 101;
			4611: Pixel = 103;
			4612: Pixel = 110;
			4613: Pixel = 115;
			4614: Pixel = 111;
			4615: Pixel = 95;
			4616: Pixel = 195;
			4617: Pixel = 197;
			4618: Pixel = 102;
			4619: Pixel = 110;
			4620: Pixel = 115;
			4621: Pixel = 118;
			4622: Pixel = 125;
			4623: Pixel = 114;
			4624: Pixel = 117;
			4625: Pixel = 85;
			4626: Pixel = 50;
			4627: Pixel = 66;
			4628: Pixel = 42;
			4629: Pixel = 47;
			4630: Pixel = 59;
			4631: Pixel = 76;
			4632: Pixel = 68;
			4633: Pixel = 56;
			4634: Pixel = 68;
			4635: Pixel = 104;
			4636: Pixel = 57;
			4637: Pixel = 29;
			4638: Pixel = 61;
			4639: Pixel = 126;
			4640: Pixel = 139;
			4641: Pixel = 157;
			4642: Pixel = 157;
			4643: Pixel = 184;
			4644: Pixel = 188;
			4645: Pixel = 173;
			4646: Pixel = 159;
			4647: Pixel = 174;
			4648: Pixel = 171;
			4649: Pixel = 163;
			4650: Pixel = 180;
			4651: Pixel = 193;
			4652: Pixel = 197;
			4653: Pixel = 201;
			4654: Pixel = 200;
			4655: Pixel = 205;
			4656: Pixel = 207;
			4657: Pixel = 176;
			4658: Pixel = 101;
			4659: Pixel = 47;
			4660: Pixel = 53;
			4661: Pixel = 101;
			4662: Pixel = 166;
			4663: Pixel = 83;
			4664: Pixel = 40;
			4665: Pixel = 50;
			4666: Pixel = 52;
			4667: Pixel = 55;
			4668: Pixel = 62;
			4669: Pixel = 55;
			4670: Pixel = 44;
			4671: Pixel = 50;
			4672: Pixel = 45;
			4673: Pixel = 88;
			4674: Pixel = 139;
			4675: Pixel = 135;
			4676: Pixel = 153;
			4677: Pixel = 151;
			4678: Pixel = 157;
			4679: Pixel = 162;
			4680: Pixel = 164;
			4681: Pixel = 162;
			4682: Pixel = 161;
			4683: Pixel = 161;
			4684: Pixel = 163;
			4685: Pixel = 160;
			4686: Pixel = 159;
			4687: Pixel = 157;
			4688: Pixel = 158;
			4689: Pixel = 157;
			4690: Pixel = 154;
			4691: Pixel = 151;
			4692: Pixel = 103;
			4693: Pixel = 104;
			4694: Pixel = 102;
			4695: Pixel = 100;
			4696: Pixel = 92;
			4697: Pixel = 110;
			4698: Pixel = 147;
			4699: Pixel = 166;
			4700: Pixel = 172;
			4701: Pixel = 173;
			4702: Pixel = 173;
			4703: Pixel = 156;
			4704: Pixel = 116;
			4705: Pixel = 75;
			4706: Pixel = 80;
			4707: Pixel = 92;
			4708: Pixel = 99;
			4709: Pixel = 103;
			4710: Pixel = 103;
			4711: Pixel = 101;
			4712: Pixel = 98;
			4713: Pixel = 107;
			4714: Pixel = 128;
			4715: Pixel = 113;
			4716: Pixel = 116;
			4717: Pixel = 97;
			4718: Pixel = 163;
			4719: Pixel = 184;
			4720: Pixel = 106;
			4721: Pixel = 115;
			4722: Pixel = 111;
			4723: Pixel = 131;
			4724: Pixel = 121;
			4725: Pixel = 90;
			4726: Pixel = 69;
			4727: Pixel = 55;
			4728: Pixel = 71;
			4729: Pixel = 57;
			4730: Pixel = 51;
			4731: Pixel = 55;
			4732: Pixel = 48;
			4733: Pixel = 57;
			4734: Pixel = 60;
			4735: Pixel = 86;
			4736: Pixel = 73;
			4737: Pixel = 85;
			4738: Pixel = 29;
			4739: Pixel = 48;
			4740: Pixel = 128;
			4741: Pixel = 145;
			4742: Pixel = 178;
			4743: Pixel = 158;
			4744: Pixel = 154;
			4745: Pixel = 179;
			4746: Pixel = 184;
			4747: Pixel = 169;
			4748: Pixel = 170;
			4749: Pixel = 161;
			4750: Pixel = 158;
			4751: Pixel = 174;
			4752: Pixel = 187;
			4753: Pixel = 194;
			4754: Pixel = 199;
			4755: Pixel = 201;
			4756: Pixel = 204;
			4757: Pixel = 208;
			4758: Pixel = 211;
			4759: Pixel = 194;
			4760: Pixel = 121;
			4761: Pixel = 55;
			4762: Pixel = 39;
			4763: Pixel = 74;
			4764: Pixel = 162;
			4765: Pixel = 94;
			4766: Pixel = 45;
			4767: Pixel = 54;
			4768: Pixel = 56;
			4769: Pixel = 58;
			4770: Pixel = 63;
			4771: Pixel = 49;
			4772: Pixel = 46;
			4773: Pixel = 53;
			4774: Pixel = 45;
			4775: Pixel = 116;
			4776: Pixel = 138;
			4777: Pixel = 147;
			4778: Pixel = 159;
			4779: Pixel = 151;
			4780: Pixel = 149;
			4781: Pixel = 150;
			4782: Pixel = 151;
			4783: Pixel = 155;
			4784: Pixel = 158;
			4785: Pixel = 159;
			4786: Pixel = 161;
			4787: Pixel = 161;
			4788: Pixel = 159;
			4789: Pixel = 158;
			4790: Pixel = 156;
			4791: Pixel = 156;
			4792: Pixel = 154;
			4793: Pixel = 151;
			4794: Pixel = 106;
			4795: Pixel = 103;
			4796: Pixel = 99;
			4797: Pixel = 97;
			4798: Pixel = 91;
			4799: Pixel = 109;
			4800: Pixel = 145;
			4801: Pixel = 166;
			4802: Pixel = 173;
			4803: Pixel = 174;
			4804: Pixel = 173;
			4805: Pixel = 156;
			4806: Pixel = 115;
			4807: Pixel = 78;
			4808: Pixel = 86;
			4809: Pixel = 96;
			4810: Pixel = 100;
			4811: Pixel = 102;
			4812: Pixel = 102;
			4813: Pixel = 101;
			4814: Pixel = 99;
			4815: Pixel = 112;
			4816: Pixel = 117;
			4817: Pixel = 116;
			4818: Pixel = 119;
			4819: Pixel = 114;
			4820: Pixel = 123;
			4821: Pixel = 184;
			4822: Pixel = 113;
			4823: Pixel = 117;
			4824: Pixel = 127;
			4825: Pixel = 131;
			4826: Pixel = 115;
			4827: Pixel = 75;
			4828: Pixel = 64;
			4829: Pixel = 41;
			4830: Pixel = 58;
			4831: Pixel = 66;
			4832: Pixel = 53;
			4833: Pixel = 55;
			4834: Pixel = 51;
			4835: Pixel = 55;
			4836: Pixel = 52;
			4837: Pixel = 86;
			4838: Pixel = 72;
			4839: Pixel = 98;
			4840: Pixel = 47;
			4841: Pixel = 115;
			4842: Pixel = 142;
			4843: Pixel = 175;
			4844: Pixel = 184;
			4845: Pixel = 169;
			4846: Pixel = 152;
			4847: Pixel = 188;
			4848: Pixel = 182;
			4849: Pixel = 164;
			4850: Pixel = 157;
			4851: Pixel = 156;
			4852: Pixel = 169;
			4853: Pixel = 176;
			4854: Pixel = 191;
			4855: Pixel = 195;
			4856: Pixel = 199;
			4857: Pixel = 203;
			4858: Pixel = 205;
			4859: Pixel = 209;
			4860: Pixel = 212;
			4861: Pixel = 204;
			4862: Pixel = 138;
			4863: Pixel = 66;
			4864: Pixel = 36;
			4865: Pixel = 57;
			4866: Pixel = 150;
			4867: Pixel = 107;
			4868: Pixel = 45;
			4869: Pixel = 55;
			4870: Pixel = 57;
			4871: Pixel = 60;
			4872: Pixel = 62;
			4873: Pixel = 48;
			4874: Pixel = 51;
			4875: Pixel = 47;
			4876: Pixel = 64;
			4877: Pixel = 139;
			4878: Pixel = 136;
			4879: Pixel = 160;
			4880: Pixel = 164;
			4881: Pixel = 158;
			4882: Pixel = 154;
			4883: Pixel = 151;
			4884: Pixel = 149;
			4885: Pixel = 150;
			4886: Pixel = 147;
			4887: Pixel = 148;
			4888: Pixel = 152;
			4889: Pixel = 156;
			4890: Pixel = 157;
			4891: Pixel = 156;
			4892: Pixel = 154;
			4893: Pixel = 153;
			4894: Pixel = 153;
			4895: Pixel = 150;
			4896: Pixel = 103;
			4897: Pixel = 102;
			4898: Pixel = 99;
			4899: Pixel = 97;
			4900: Pixel = 89;
			4901: Pixel = 108;
			4902: Pixel = 146;
			4903: Pixel = 167;
			4904: Pixel = 174;
			4905: Pixel = 175;
			4906: Pixel = 172;
			4907: Pixel = 157;
			4908: Pixel = 114;
			4909: Pixel = 76;
			4910: Pixel = 86;
			4911: Pixel = 95;
			4912: Pixel = 99;
			4913: Pixel = 101;
			4914: Pixel = 104;
			4915: Pixel = 103;
			4916: Pixel = 103;
			4917: Pixel = 108;
			4918: Pixel = 116;
			4919: Pixel = 116;
			4920: Pixel = 117;
			4921: Pixel = 114;
			4922: Pixel = 117;
			4923: Pixel = 133;
			4924: Pixel = 118;
			4925: Pixel = 131;
			4926: Pixel = 133;
			4927: Pixel = 121;
			4928: Pixel = 70;
			4929: Pixel = 47;
			4930: Pixel = 71;
			4931: Pixel = 54;
			4932: Pixel = 46;
			4933: Pixel = 63;
			4934: Pixel = 70;
			4935: Pixel = 51;
			4936: Pixel = 48;
			4937: Pixel = 65;
			4938: Pixel = 52;
			4939: Pixel = 64;
			4940: Pixel = 52;
			4941: Pixel = 49;
			4942: Pixel = 117;
			4943: Pixel = 134;
			4944: Pixel = 159;
			4945: Pixel = 168;
			4946: Pixel = 188;
			4947: Pixel = 176;
			4948: Pixel = 153;
			4949: Pixel = 188;
			4950: Pixel = 162;
			4951: Pixel = 155;
			4952: Pixel = 157;
			4953: Pixel = 168;
			4954: Pixel = 173;
			4955: Pixel = 177;
			4956: Pixel = 187;
			4957: Pixel = 196;
			4958: Pixel = 198;
			4959: Pixel = 200;
			4960: Pixel = 204;
			4961: Pixel = 208;
			4962: Pixel = 212;
			4963: Pixel = 211;
			4964: Pixel = 157;
			4965: Pixel = 86;
			4966: Pixel = 44;
			4967: Pixel = 45;
			4968: Pixel = 137;
			4969: Pixel = 117;
			4970: Pixel = 42;
			4971: Pixel = 55;
			4972: Pixel = 59;
			4973: Pixel = 61;
			4974: Pixel = 56;
			4975: Pixel = 48;
			4976: Pixel = 53;
			4977: Pixel = 42;
			4978: Pixel = 99;
			4979: Pixel = 143;
			4980: Pixel = 141;
			4981: Pixel = 164;
			4982: Pixel = 162;
			4983: Pixel = 161;
			4984: Pixel = 161;
			4985: Pixel = 161;
			4986: Pixel = 158;
			4987: Pixel = 155;
			4988: Pixel = 150;
			4989: Pixel = 144;
			4990: Pixel = 146;
			4991: Pixel = 145;
			4992: Pixel = 145;
			4993: Pixel = 147;
			4994: Pixel = 150;
			4995: Pixel = 153;
			4996: Pixel = 154;
			4997: Pixel = 151;
			4998: Pixel = 102;
			4999: Pixel = 101;
			5000: Pixel = 98;
			5001: Pixel = 98;
			5002: Pixel = 90;
			5003: Pixel = 108;
			5004: Pixel = 147;
			5005: Pixel = 167;
			5006: Pixel = 173;
			5007: Pixel = 175;
			5008: Pixel = 174;
			5009: Pixel = 156;
			5010: Pixel = 114;
			5011: Pixel = 76;
			5012: Pixel = 83;
			5013: Pixel = 95;
			5014: Pixel = 101;
			5015: Pixel = 102;
			5016: Pixel = 103;
			5017: Pixel = 102;
			5018: Pixel = 103;
			5019: Pixel = 108;
			5020: Pixel = 115;
			5021: Pixel = 118;
			5022: Pixel = 116;
			5023: Pixel = 121;
			5024: Pixel = 131;
			5025: Pixel = 122;
			5026: Pixel = 129;
			5027: Pixel = 123;
			5028: Pixel = 131;
			5029: Pixel = 95;
			5030: Pixel = 68;
			5031: Pixel = 51;
			5032: Pixel = 74;
			5033: Pixel = 56;
			5034: Pixel = 49;
			5035: Pixel = 80;
			5036: Pixel = 67;
			5037: Pixel = 41;
			5038: Pixel = 55;
			5039: Pixel = 57;
			5040: Pixel = 65;
			5041: Pixel = 69;
			5042: Pixel = 49;
			5043: Pixel = 70;
			5044: Pixel = 120;
			5045: Pixel = 160;
			5046: Pixel = 168;
			5047: Pixel = 161;
			5048: Pixel = 184;
			5049: Pixel = 187;
			5050: Pixel = 178;
			5051: Pixel = 148;
			5052: Pixel = 151;
			5053: Pixel = 167;
			5054: Pixel = 170;
			5055: Pixel = 174;
			5056: Pixel = 176;
			5057: Pixel = 176;
			5058: Pixel = 182;
			5059: Pixel = 193;
			5060: Pixel = 196;
			5061: Pixel = 196;
			5062: Pixel = 201;
			5063: Pixel = 204;
			5064: Pixel = 209;
			5065: Pixel = 214;
			5066: Pixel = 177;
			5067: Pixel = 90;
			5068: Pixel = 44;
			5069: Pixel = 39;
			5070: Pixel = 119;
			5071: Pixel = 132;
			5072: Pixel = 52;
			5073: Pixel = 61;
			5074: Pixel = 60;
			5075: Pixel = 65;
			5076: Pixel = 51;
			5077: Pixel = 52;
			5078: Pixel = 50;
			5079: Pixel = 54;
			5080: Pixel = 126;
			5081: Pixel = 135;
			5082: Pixel = 149;
			5083: Pixel = 164;
			5084: Pixel = 161;
			5085: Pixel = 160;
			5086: Pixel = 161;
			5087: Pixel = 165;
			5088: Pixel = 166;
			5089: Pixel = 160;
			5090: Pixel = 156;
			5091: Pixel = 150;
			5092: Pixel = 148;
			5093: Pixel = 144;
			5094: Pixel = 142;
			5095: Pixel = 142;
			5096: Pixel = 142;
			5097: Pixel = 145;
			5098: Pixel = 147;
			5099: Pixel = 150;
			5100: Pixel = 101;
			5101: Pixel = 99;
			5102: Pixel = 99;
			5103: Pixel = 99;
			5104: Pixel = 91;
			5105: Pixel = 107;
			5106: Pixel = 146;
			5107: Pixel = 166;
			5108: Pixel = 174;
			5109: Pixel = 176;
			5110: Pixel = 174;
			5111: Pixel = 157;
			5112: Pixel = 115;
			5113: Pixel = 76;
			5114: Pixel = 84;
			5115: Pixel = 93;
			5116: Pixel = 101;
			5117: Pixel = 103;
			5118: Pixel = 102;
			5119: Pixel = 101;
			5120: Pixel = 102;
			5121: Pixel = 109;
			5122: Pixel = 117;
			5123: Pixel = 118;
			5124: Pixel = 121;
			5125: Pixel = 165;
			5126: Pixel = 86;
			5127: Pixel = 47;
			5128: Pixel = 133;
			5129: Pixel = 143;
			5130: Pixel = 99;
			5131: Pixel = 68;
			5132: Pixel = 81;
			5133: Pixel = 47;
			5134: Pixel = 95;
			5135: Pixel = 41;
			5136: Pixel = 55;
			5137: Pixel = 62;
			5138: Pixel = 45;
			5139: Pixel = 46;
			5140: Pixel = 59;
			5141: Pixel = 60;
			5142: Pixel = 73;
			5143: Pixel = 56;
			5144: Pixel = 55;
			5145: Pixel = 120;
			5146: Pixel = 150;
			5147: Pixel = 182;
			5148: Pixel = 176;
			5149: Pixel = 156;
			5150: Pixel = 192;
			5151: Pixel = 190;
			5152: Pixel = 130;
			5153: Pixel = 102;
			5154: Pixel = 109;
			5155: Pixel = 107;
			5156: Pixel = 131;
			5157: Pixel = 168;
			5158: Pixel = 183;
			5159: Pixel = 176;
			5160: Pixel = 176;
			5161: Pixel = 187;
			5162: Pixel = 194;
			5163: Pixel = 190;
			5164: Pixel = 196;
			5165: Pixel = 203;
			5166: Pixel = 210;
			5167: Pixel = 191;
			5168: Pixel = 139;
			5169: Pixel = 65;
			5170: Pixel = 40;
			5171: Pixel = 38;
			5172: Pixel = 101;
			5173: Pixel = 147;
			5174: Pixel = 57;
			5175: Pixel = 62;
			5176: Pixel = 63;
			5177: Pixel = 63;
			5178: Pixel = 48;
			5179: Pixel = 53;
			5180: Pixel = 46;
			5181: Pixel = 74;
			5182: Pixel = 138;
			5183: Pixel = 133;
			5184: Pixel = 158;
			5185: Pixel = 160;
			5186: Pixel = 158;
			5187: Pixel = 158;
			5188: Pixel = 158;
			5189: Pixel = 159;
			5190: Pixel = 161;
			5191: Pixel = 161;
			5192: Pixel = 155;
			5193: Pixel = 155;
			5194: Pixel = 153;
			5195: Pixel = 150;
			5196: Pixel = 149;
			5197: Pixel = 147;
			5198: Pixel = 141;
			5199: Pixel = 140;
			5200: Pixel = 139;
			5201: Pixel = 137;
			5202: Pixel = 102;
			5203: Pixel = 102;
			5204: Pixel = 102;
			5205: Pixel = 100;
			5206: Pixel = 91;
			5207: Pixel = 105;
			5208: Pixel = 145;
			5209: Pixel = 166;
			5210: Pixel = 174;
			5211: Pixel = 176;
			5212: Pixel = 175;
			5213: Pixel = 158;
			5214: Pixel = 115;
			5215: Pixel = 77;
			5216: Pixel = 85;
			5217: Pixel = 94;
			5218: Pixel = 101;
			5219: Pixel = 102;
			5220: Pixel = 100;
			5221: Pixel = 100;
			5222: Pixel = 102;
			5223: Pixel = 108;
			5224: Pixel = 110;
			5225: Pixel = 120;
			5226: Pixel = 139;
			5227: Pixel = 149;
			5228: Pixel = 66;
			5229: Pixel = 44;
			5230: Pixel = 137;
			5231: Pixel = 111;
			5232: Pixel = 62;
			5233: Pixel = 77;
			5234: Pixel = 67;
			5235: Pixel = 66;
			5236: Pixel = 94;
			5237: Pixel = 45;
			5238: Pixel = 58;
			5239: Pixel = 61;
			5240: Pixel = 67;
			5241: Pixel = 40;
			5242: Pixel = 44;
			5243: Pixel = 80;
			5244: Pixel = 72;
			5245: Pixel = 38;
			5246: Pixel = 108;
			5247: Pixel = 147;
			5248: Pixel = 173;
			5249: Pixel = 190;
			5250: Pixel = 166;
			5251: Pixel = 177;
			5252: Pixel = 188;
			5253: Pixel = 135;
			5254: Pixel = 140;
			5255: Pixel = 148;
			5256: Pixel = 148;
			5257: Pixel = 104;
			5258: Pixel = 75;
			5259: Pixel = 85;
			5260: Pixel = 143;
			5261: Pixel = 172;
			5262: Pixel = 170;
			5263: Pixel = 183;
			5264: Pixel = 191;
			5265: Pixel = 188;
			5266: Pixel = 191;
			5267: Pixel = 180;
			5268: Pixel = 140;
			5269: Pixel = 108;
			5270: Pixel = 103;
			5271: Pixel = 90;
			5272: Pixel = 53;
			5273: Pixel = 39;
			5274: Pixel = 84;
			5275: Pixel = 156;
			5276: Pixel = 61;
			5277: Pixel = 61;
			5278: Pixel = 66;
			5279: Pixel = 55;
			5280: Pixel = 49;
			5281: Pixel = 54;
			5282: Pixel = 49;
			5283: Pixel = 96;
			5284: Pixel = 137;
			5285: Pixel = 139;
			5286: Pixel = 163;
			5287: Pixel = 159;
			5288: Pixel = 157;
			5289: Pixel = 157;
			5290: Pixel = 155;
			5291: Pixel = 155;
			5292: Pixel = 157;
			5293: Pixel = 158;
			5294: Pixel = 155;
			5295: Pixel = 153;
			5296: Pixel = 154;
			5297: Pixel = 155;
			5298: Pixel = 155;
			5299: Pixel = 152;
			5300: Pixel = 147;
			5301: Pixel = 144;
			5302: Pixel = 138;
			5303: Pixel = 132;
			5304: Pixel = 101;
			5305: Pixel = 103;
			5306: Pixel = 102;
			5307: Pixel = 99;
			5308: Pixel = 86;
			5309: Pixel = 105;
			5310: Pixel = 145;
			5311: Pixel = 166;
			5312: Pixel = 175;
			5313: Pixel = 175;
			5314: Pixel = 175;
			5315: Pixel = 160;
			5316: Pixel = 118;
			5317: Pixel = 76;
			5318: Pixel = 84;
			5319: Pixel = 95;
			5320: Pixel = 102;
			5321: Pixel = 102;
			5322: Pixel = 100;
			5323: Pixel = 99;
			5324: Pixel = 100;
			5325: Pixel = 99;
			5326: Pixel = 115;
			5327: Pixel = 140;
			5328: Pixel = 154;
			5329: Pixel = 154;
			5330: Pixel = 152;
			5331: Pixel = 122;
			5332: Pixel = 86;
			5333: Pixel = 65;
			5334: Pixel = 69;
			5335: Pixel = 92;
			5336: Pixel = 75;
			5337: Pixel = 76;
			5338: Pixel = 59;
			5339: Pixel = 65;
			5340: Pixel = 57;
			5341: Pixel = 40;
			5342: Pixel = 86;
			5343: Pixel = 48;
			5344: Pixel = 38;
			5345: Pixel = 50;
			5346: Pixel = 43;
			5347: Pixel = 71;
			5348: Pixel = 141;
			5349: Pixel = 172;
			5350: Pixel = 184;
			5351: Pixel = 193;
			5352: Pixel = 179;
			5353: Pixel = 173;
			5354: Pixel = 101;
			5355: Pixel = 91;
			5356: Pixel = 93;
			5357: Pixel = 74;
			5358: Pixel = 89;
			5359: Pixel = 82;
			5360: Pixel = 112;
			5361: Pixel = 110;
			5362: Pixel = 114;
			5363: Pixel = 151;
			5364: Pixel = 160;
			5365: Pixel = 179;
			5366: Pixel = 194;
			5367: Pixel = 194;
			5368: Pixel = 182;
			5369: Pixel = 123;
			5370: Pixel = 80;
			5371: Pixel = 71;
			5372: Pixel = 84;
			5373: Pixel = 79;
			5374: Pixel = 62;
			5375: Pixel = 38;
			5376: Pixel = 81;
			5377: Pixel = 155;
			5378: Pixel = 72;
			5379: Pixel = 57;
			5380: Pixel = 65;
			5381: Pixel = 51;
			5382: Pixel = 50;
			5383: Pixel = 51;
			5384: Pixel = 51;
			5385: Pixel = 121;
			5386: Pixel = 134;
			5387: Pixel = 149;
			5388: Pixel = 161;
			5389: Pixel = 157;
			5390: Pixel = 156;
			5391: Pixel = 156;
			5392: Pixel = 155;
			5393: Pixel = 154;
			5394: Pixel = 156;
			5395: Pixel = 157;
			5396: Pixel = 154;
			5397: Pixel = 152;
			5398: Pixel = 153;
			5399: Pixel = 154;
			5400: Pixel = 156;
			5401: Pixel = 154;
			5402: Pixel = 149;
			5403: Pixel = 148;
			5404: Pixel = 141;
			5405: Pixel = 135;
			5406: Pixel = 98;
			5407: Pixel = 97;
			5408: Pixel = 96;
			5409: Pixel = 94;
			5410: Pixel = 82;
			5411: Pixel = 99;
			5412: Pixel = 144;
			5413: Pixel = 167;
			5414: Pixel = 176;
			5415: Pixel = 177;
			5416: Pixel = 173;
			5417: Pixel = 157;
			5418: Pixel = 118;
			5419: Pixel = 74;
			5420: Pixel = 81;
			5421: Pixel = 90;
			5422: Pixel = 98;
			5423: Pixel = 100;
			5424: Pixel = 97;
			5425: Pixel = 97;
			5426: Pixel = 87;
			5427: Pixel = 135;
			5428: Pixel = 176;
			5429: Pixel = 141;
			5430: Pixel = 152;
			5431: Pixel = 150;
			5432: Pixel = 110;
			5433: Pixel = 72;
			5434: Pixel = 39;
			5435: Pixel = 80;
			5436: Pixel = 92;
			5437: Pixel = 82;
			5438: Pixel = 92;
			5439: Pixel = 81;
			5440: Pixel = 47;
			5441: Pixel = 64;
			5442: Pixel = 73;
			5443: Pixel = 36;
			5444: Pixel = 56;
			5445: Pixel = 94;
			5446: Pixel = 55;
			5447: Pixel = 38;
			5448: Pixel = 40;
			5449: Pixel = 122;
			5450: Pixel = 165;
			5451: Pixel = 175;
			5452: Pixel = 192;
			5453: Pixel = 198;
			5454: Pixel = 171;
			5455: Pixel = 78;
			5456: Pixel = 51;
			5457: Pixel = 50;
			5458: Pixel = 42;
			5459: Pixel = 49;
			5460: Pixel = 86;
			5461: Pixel = 43;
			5462: Pixel = 53;
			5463: Pixel = 127;
			5464: Pixel = 132;
			5465: Pixel = 139;
			5466: Pixel = 153;
			5467: Pixel = 178;
			5468: Pixel = 203;
			5469: Pixel = 198;
			5470: Pixel = 105;
			5471: Pixel = 54;
			5472: Pixel = 69;
			5473: Pixel = 59;
			5474: Pixel = 45;
			5475: Pixel = 58;
			5476: Pixel = 51;
			5477: Pixel = 39;
			5478: Pixel = 75;
			5479: Pixel = 154;
			5480: Pixel = 81;
			5481: Pixel = 62;
			5482: Pixel = 60;
			5483: Pixel = 47;
			5484: Pixel = 51;
			5485: Pixel = 48;
			5486: Pixel = 59;
			5487: Pixel = 137;
			5488: Pixel = 138;
			5489: Pixel = 157;
			5490: Pixel = 158;
			5491: Pixel = 155;
			5492: Pixel = 153;
			5493: Pixel = 154;
			5494: Pixel = 155;
			5495: Pixel = 154;
			5496: Pixel = 155;
			5497: Pixel = 155;
			5498: Pixel = 153;
			5499: Pixel = 153;
			5500: Pixel = 153;
			5501: Pixel = 151;
			5502: Pixel = 153;
			5503: Pixel = 148;
			5504: Pixel = 144;
			5505: Pixel = 142;
			5506: Pixel = 141;
			5507: Pixel = 136;
			5508: Pixel = 97;
			5509: Pixel = 95;
			5510: Pixel = 93;
			5511: Pixel = 89;
			5512: Pixel = 76;
			5513: Pixel = 95;
			5514: Pixel = 143;
			5515: Pixel = 169;
			5516: Pixel = 176;
			5517: Pixel = 177;
			5518: Pixel = 176;
			5519: Pixel = 156;
			5520: Pixel = 116;
			5521: Pixel = 74;
			5522: Pixel = 84;
			5523: Pixel = 95;
			5524: Pixel = 98;
			5525: Pixel = 97;
			5526: Pixel = 99;
			5527: Pixel = 99;
			5528: Pixel = 80;
			5529: Pixel = 156;
			5530: Pixel = 167;
			5531: Pixel = 138;
			5532: Pixel = 150;
			5533: Pixel = 129;
			5534: Pixel = 69;
			5535: Pixel = 41;
			5536: Pixel = 78;
			5537: Pixel = 72;
			5538: Pixel = 57;
			5539: Pixel = 63;
			5540: Pixel = 111;
			5541: Pixel = 70;
			5542: Pixel = 43;
			5543: Pixel = 44;
			5544: Pixel = 80;
			5545: Pixel = 55;
			5546: Pixel = 38;
			5547: Pixel = 55;
			5548: Pixel = 62;
			5549: Pixel = 40;
			5550: Pixel = 84;
			5551: Pixel = 147;
			5552: Pixel = 174;
			5553: Pixel = 179;
			5554: Pixel = 203;
			5555: Pixel = 187;
			5556: Pixel = 97;
			5557: Pixel = 53;
			5558: Pixel = 52;
			5559: Pixel = 75;
			5560: Pixel = 57;
			5561: Pixel = 61;
			5562: Pixel = 180;
			5563: Pixel = 162;
			5564: Pixel = 67;
			5565: Pixel = 102;
			5566: Pixel = 123;
			5567: Pixel = 134;
			5568: Pixel = 148;
			5569: Pixel = 180;
			5570: Pixel = 220;
			5571: Pixel = 135;
			5572: Pixel = 43;
			5573: Pixel = 53;
			5574: Pixel = 112;
			5575: Pixel = 133;
			5576: Pixel = 47;
			5577: Pixel = 50;
			5578: Pixel = 48;
			5579: Pixel = 45;
			5580: Pixel = 72;
			5581: Pixel = 152;
			5582: Pixel = 88;
			5583: Pixel = 69;
			5584: Pixel = 57;
			5585: Pixel = 48;
			5586: Pixel = 52;
			5587: Pixel = 43;
			5588: Pixel = 91;
			5589: Pixel = 143;
			5590: Pixel = 144;
			5591: Pixel = 159;
			5592: Pixel = 156;
			5593: Pixel = 154;
			5594: Pixel = 152;
			5595: Pixel = 152;
			5596: Pixel = 152;
			5597: Pixel = 153;
			5598: Pixel = 152;
			5599: Pixel = 153;
			5600: Pixel = 152;
			5601: Pixel = 152;
			5602: Pixel = 150;
			5603: Pixel = 148;
			5604: Pixel = 147;
			5605: Pixel = 143;
			5606: Pixel = 139;
			5607: Pixel = 133;
			5608: Pixel = 130;
			5609: Pixel = 131;
			5610: Pixel = 99;
			5611: Pixel = 97;
			5612: Pixel = 96;
			5613: Pixel = 90;
			5614: Pixel = 74;
			5615: Pixel = 93;
			5616: Pixel = 143;
			5617: Pixel = 168;
			5618: Pixel = 177;
			5619: Pixel = 179;
			5620: Pixel = 178;
			5621: Pixel = 158;
			5622: Pixel = 117;
			5623: Pixel = 80;
			5624: Pixel = 87;
			5625: Pixel = 100;
			5626: Pixel = 104;
			5627: Pixel = 102;
			5628: Pixel = 106;
			5629: Pixel = 91;
			5630: Pixel = 55;
			5631: Pixel = 104;
			5632: Pixel = 162;
			5633: Pixel = 214;
			5634: Pixel = 118;
			5635: Pixel = 47;
			5636: Pixel = 43;
			5637: Pixel = 84;
			5638: Pixel = 64;
			5639: Pixel = 63;
			5640: Pixel = 68;
			5641: Pixel = 86;
			5642: Pixel = 113;
			5643: Pixel = 72;
			5644: Pixel = 41;
			5645: Pixel = 44;
			5646: Pixel = 61;
			5647: Pixel = 60;
			5648: Pixel = 44;
			5649: Pixel = 46;
			5650: Pixel = 33;
			5651: Pixel = 55;
			5652: Pixel = 112;
			5653: Pixel = 156;
			5654: Pixel = 171;
			5655: Pixel = 198;
			5656: Pixel = 192;
			5657: Pixel = 122;
			5658: Pixel = 117;
			5659: Pixel = 106;
			5660: Pixel = 66;
			5661: Pixel = 107;
			5662: Pixel = 89;
			5663: Pixel = 113;
			5664: Pixel = 208;
			5665: Pixel = 200;
			5666: Pixel = 122;
			5667: Pixel = 111;
			5668: Pixel = 116;
			5669: Pixel = 128;
			5670: Pixel = 147;
			5671: Pixel = 197;
			5672: Pixel = 204;
			5673: Pixel = 108;
			5674: Pixel = 102;
			5675: Pixel = 85;
			5676: Pixel = 139;
			5677: Pixel = 152;
			5678: Pixel = 54;
			5679: Pixel = 45;
			5680: Pixel = 45;
			5681: Pixel = 50;
			5682: Pixel = 71;
			5683: Pixel = 152;
			5684: Pixel = 95;
			5685: Pixel = 74;
			5686: Pixel = 51;
			5687: Pixel = 50;
			5688: Pixel = 52;
			5689: Pixel = 44;
			5690: Pixel = 115;
			5691: Pixel = 142;
			5692: Pixel = 150;
			5693: Pixel = 158;
			5694: Pixel = 155;
			5695: Pixel = 153;
			5696: Pixel = 151;
			5697: Pixel = 152;
			5698: Pixel = 152;
			5699: Pixel = 153;
			5700: Pixel = 152;
			5701: Pixel = 152;
			5702: Pixel = 151;
			5703: Pixel = 149;
			5704: Pixel = 147;
			5705: Pixel = 145;
			5706: Pixel = 142;
			5707: Pixel = 137;
			5708: Pixel = 130;
			5709: Pixel = 130;
			5710: Pixel = 142;
			5711: Pixel = 161;
			5712: Pixel = 102;
			5713: Pixel = 100;
			5714: Pixel = 96;
			5715: Pixel = 89;
			5716: Pixel = 75;
			5717: Pixel = 92;
			5718: Pixel = 144;
			5719: Pixel = 167;
			5720: Pixel = 178;
			5721: Pixel = 180;
			5722: Pixel = 179;
			5723: Pixel = 160;
			5724: Pixel = 119;
			5725: Pixel = 84;
			5726: Pixel = 92;
			5727: Pixel = 104;
			5728: Pixel = 108;
			5729: Pixel = 118;
			5730: Pixel = 67;
			5731: Pixel = 63;
			5732: Pixel = 128;
			5733: Pixel = 157;
			5734: Pixel = 181;
			5735: Pixel = 119;
			5736: Pixel = 60;
			5737: Pixel = 70;
			5738: Pixel = 84;
			5739: Pixel = 82;
			5740: Pixel = 42;
			5741: Pixel = 78;
			5742: Pixel = 78;
			5743: Pixel = 98;
			5744: Pixel = 118;
			5745: Pixel = 99;
			5746: Pixel = 54;
			5747: Pixel = 42;
			5748: Pixel = 44;
			5749: Pixel = 49;
			5750: Pixel = 50;
			5751: Pixel = 47;
			5752: Pixel = 32;
			5753: Pixel = 94;
			5754: Pixel = 151;
			5755: Pixel = 174;
			5756: Pixel = 194;
			5757: Pixel = 193;
			5758: Pixel = 119;
			5759: Pixel = 121;
			5760: Pixel = 136;
			5761: Pixel = 146;
			5762: Pixel = 121;
			5763: Pixel = 113;
			5764: Pixel = 123;
			5765: Pixel = 153;
			5766: Pixel = 168;
			5767: Pixel = 168;
			5768: Pixel = 151;
			5769: Pixel = 128;
			5770: Pixel = 122;
			5771: Pixel = 127;
			5772: Pixel = 144;
			5773: Pixel = 202;
			5774: Pixel = 205;
			5775: Pixel = 131;
			5776: Pixel = 134;
			5777: Pixel = 136;
			5778: Pixel = 152;
			5779: Pixel = 96;
			5780: Pixel = 61;
			5781: Pixel = 60;
			5782: Pixel = 49;
			5783: Pixel = 59;
			5784: Pixel = 65;
			5785: Pixel = 153;
			5786: Pixel = 105;
			5787: Pixel = 71;
			5788: Pixel = 48;
			5789: Pixel = 48;
			5790: Pixel = 51;
			5791: Pixel = 64;
			5792: Pixel = 131;
			5793: Pixel = 140;
			5794: Pixel = 155;
			5795: Pixel = 156;
			5796: Pixel = 153;
			5797: Pixel = 151;
			5798: Pixel = 149;
			5799: Pixel = 156;
			5800: Pixel = 156;
			5801: Pixel = 151;
			5802: Pixel = 154;
			5803: Pixel = 151;
			5804: Pixel = 148;
			5805: Pixel = 145;
			5806: Pixel = 142;
			5807: Pixel = 139;
			5808: Pixel = 136;
			5809: Pixel = 133;
			5810: Pixel = 145;
			5811: Pixel = 167;
			5812: Pixel = 180;
			5813: Pixel = 187;
			5814: Pixel = 102;
			5815: Pixel = 101;
			5816: Pixel = 93;
			5817: Pixel = 86;
			5818: Pixel = 72;
			5819: Pixel = 89;
			5820: Pixel = 143;
			5821: Pixel = 168;
			5822: Pixel = 177;
			5823: Pixel = 182;
			5824: Pixel = 182;
			5825: Pixel = 163;
			5826: Pixel = 122;
			5827: Pixel = 81;
			5828: Pixel = 91;
			5829: Pixel = 104;
			5830: Pixel = 109;
			5831: Pixel = 116;
			5832: Pixel = 110;
			5833: Pixel = 140;
			5834: Pixel = 144;
			5835: Pixel = 98;
			5836: Pixel = 94;
			5837: Pixel = 42;
			5838: Pixel = 43;
			5839: Pixel = 99;
			5840: Pixel = 116;
			5841: Pixel = 86;
			5842: Pixel = 47;
			5843: Pixel = 74;
			5844: Pixel = 82;
			5845: Pixel = 85;
			5846: Pixel = 120;
			5847: Pixel = 117;
			5848: Pixel = 62;
			5849: Pixel = 44;
			5850: Pixel = 47;
			5851: Pixel = 46;
			5852: Pixel = 50;
			5853: Pixel = 32;
			5854: Pixel = 62;
			5855: Pixel = 128;
			5856: Pixel = 162;
			5857: Pixel = 183;
			5858: Pixel = 199;
			5859: Pixel = 111;
			5860: Pixel = 111;
			5861: Pixel = 141;
			5862: Pixel = 145;
			5863: Pixel = 146;
			5864: Pixel = 147;
			5865: Pixel = 139;
			5866: Pixel = 125;
			5867: Pixel = 129;
			5868: Pixel = 131;
			5869: Pixel = 153;
			5870: Pixel = 158;
			5871: Pixel = 131;
			5872: Pixel = 129;
			5873: Pixel = 128;
			5874: Pixel = 138;
			5875: Pixel = 193;
			5876: Pixel = 215;
			5877: Pixel = 166;
			5878: Pixel = 140;
			5879: Pixel = 127;
			5880: Pixel = 106;
			5881: Pixel = 81;
			5882: Pixel = 92;
			5883: Pixel = 64;
			5884: Pixel = 44;
			5885: Pixel = 60;
			5886: Pixel = 60;
			5887: Pixel = 153;
			5888: Pixel = 117;
			5889: Pixel = 62;
			5890: Pixel = 47;
			5891: Pixel = 53;
			5892: Pixel = 47;
			5893: Pixel = 88;
			5894: Pixel = 138;
			5895: Pixel = 142;
			5896: Pixel = 159;
			5897: Pixel = 154;
			5898: Pixel = 152;
			5899: Pixel = 151;
			5900: Pixel = 150;
			5901: Pixel = 151;
			5902: Pixel = 151;
			5903: Pixel = 150;
			5904: Pixel = 151;
			5905: Pixel = 149;
			5906: Pixel = 145;
			5907: Pixel = 141;
			5908: Pixel = 138;
			5909: Pixel = 132;
			5910: Pixel = 140;
			5911: Pixel = 165;
			5912: Pixel = 184;
			5913: Pixel = 190;
			5914: Pixel = 189;
			5915: Pixel = 188;
			5916: Pixel = 98;
			5917: Pixel = 92;
			5918: Pixel = 86;
			5919: Pixel = 82;
			5920: Pixel = 64;
			5921: Pixel = 82;
			5922: Pixel = 141;
			5923: Pixel = 166;
			5924: Pixel = 178;
			5925: Pixel = 182;
			5926: Pixel = 181;
			5927: Pixel = 163;
			5928: Pixel = 123;
			5929: Pixel = 81;
			5930: Pixel = 90;
			5931: Pixel = 103;
			5932: Pixel = 108;
			5933: Pixel = 104;
			5934: Pixel = 135;
			5935: Pixel = 139;
			5936: Pixel = 95;
			5937: Pixel = 80;
			5938: Pixel = 67;
			5939: Pixel = 49;
			5940: Pixel = 68;
			5941: Pixel = 88;
			5942: Pixel = 101;
			5943: Pixel = 89;
			5944: Pixel = 41;
			5945: Pixel = 68;
			5946: Pixel = 80;
			5947: Pixel = 106;
			5948: Pixel = 94;
			5949: Pixel = 107;
			5950: Pixel = 56;
			5951: Pixel = 45;
			5952: Pixel = 45;
			5953: Pixel = 48;
			5954: Pixel = 49;
			5955: Pixel = 39;
			5956: Pixel = 106;
			5957: Pixel = 143;
			5958: Pixel = 181;
			5959: Pixel = 203;
			5960: Pixel = 118;
			5961: Pixel = 92;
			5962: Pixel = 128;
			5963: Pixel = 140;
			5964: Pixel = 153;
			5965: Pixel = 158;
			5966: Pixel = 160;
			5967: Pixel = 158;
			5968: Pixel = 156;
			5969: Pixel = 161;
			5970: Pixel = 168;
			5971: Pixel = 167;
			5972: Pixel = 159;
			5973: Pixel = 137;
			5974: Pixel = 137;
			5975: Pixel = 127;
			5976: Pixel = 134;
			5977: Pixel = 189;
			5978: Pixel = 216;
			5979: Pixel = 180;
			5980: Pixel = 157;
			5981: Pixel = 144;
			5982: Pixel = 130;
			5983: Pixel = 119;
			5984: Pixel = 109;
			5985: Pixel = 70;
			5986: Pixel = 46;
			5987: Pixel = 60;
			5988: Pixel = 55;
			5989: Pixel = 152;
			5990: Pixel = 122;
			5991: Pixel = 56;
			5992: Pixel = 48;
			5993: Pixel = 51;
			5994: Pixel = 42;
			5995: Pixel = 104;
			5996: Pixel = 138;
			5997: Pixel = 148;
			5998: Pixel = 157;
			5999: Pixel = 153;
			6000: Pixel = 151;
			6001: Pixel = 150;
			6002: Pixel = 151;
			6003: Pixel = 150;
			6004: Pixel = 149;
			6005: Pixel = 149;
			6006: Pixel = 147;
			6007: Pixel = 145;
			6008: Pixel = 143;
			6009: Pixel = 140;
			6010: Pixel = 131;
			6011: Pixel = 142;
			6012: Pixel = 180;
			6013: Pixel = 195;
			6014: Pixel = 193;
			6015: Pixel = 190;
			6016: Pixel = 188;
			6017: Pixel = 189;
			6018: Pixel = 93;
			6019: Pixel = 89;
			6020: Pixel = 83;
			6021: Pixel = 78;
			6022: Pixel = 61;
			6023: Pixel = 81;
			6024: Pixel = 139;
			6025: Pixel = 166;
			6026: Pixel = 177;
			6027: Pixel = 180;
			6028: Pixel = 180;
			6029: Pixel = 163;
			6030: Pixel = 122;
			6031: Pixel = 81;
			6032: Pixel = 89;
			6033: Pixel = 99;
			6034: Pixel = 113;
			6035: Pixel = 127;
			6036: Pixel = 133;
			6037: Pixel = 134;
			6038: Pixel = 115;
			6039: Pixel = 96;
			6040: Pixel = 54;
			6041: Pixel = 69;
			6042: Pixel = 97;
			6043: Pixel = 109;
			6044: Pixel = 96;
			6045: Pixel = 56;
			6046: Pixel = 36;
			6047: Pixel = 70;
			6048: Pixel = 91;
			6049: Pixel = 105;
			6050: Pixel = 113;
			6051: Pixel = 105;
			6052: Pixel = 81;
			6053: Pixel = 55;
			6054: Pixel = 46;
			6055: Pixel = 47;
			6056: Pixel = 40;
			6057: Pixel = 76;
			6058: Pixel = 126;
			6059: Pixel = 163;
			6060: Pixel = 207;
			6061: Pixel = 135;
			6062: Pixel = 65;
			6063: Pixel = 118;
			6064: Pixel = 126;
			6065: Pixel = 139;
			6066: Pixel = 151;
			6067: Pixel = 162;
			6068: Pixel = 169;
			6069: Pixel = 174;
			6070: Pixel = 172;
			6071: Pixel = 173;
			6072: Pixel = 172;
			6073: Pixel = 172;
			6074: Pixel = 155;
			6075: Pixel = 142;
			6076: Pixel = 138;
			6077: Pixel = 128;
			6078: Pixel = 130;
			6079: Pixel = 180;
			6080: Pixel = 218;
			6081: Pixel = 185;
			6082: Pixel = 164;
			6083: Pixel = 146;
			6084: Pixel = 134;
			6085: Pixel = 127;
			6086: Pixel = 117;
			6087: Pixel = 73;
			6088: Pixel = 49;
			6089: Pixel = 64;
			6090: Pixel = 48;
			6091: Pixel = 147;
			6092: Pixel = 132;
			6093: Pixel = 46;
			6094: Pixel = 49;
			6095: Pixel = 48;
			6096: Pixel = 52;
			6097: Pixel = 124;
			6098: Pixel = 138;
			6099: Pixel = 155;
			6100: Pixel = 156;
			6101: Pixel = 153;
			6102: Pixel = 151;
			6103: Pixel = 151;
			6104: Pixel = 151;
			6105: Pixel = 150;
			6106: Pixel = 147;
			6107: Pixel = 147;
			6108: Pixel = 145;
			6109: Pixel = 142;
			6110: Pixel = 140;
			6111: Pixel = 133;
			6112: Pixel = 141;
			6113: Pixel = 181;
			6114: Pixel = 198;
			6115: Pixel = 196;
			6116: Pixel = 192;
			6117: Pixel = 189;
			6118: Pixel = 189;
			6119: Pixel = 191;
			6120: Pixel = 87;
			6121: Pixel = 83;
			6122: Pixel = 79;
			6123: Pixel = 76;
			6124: Pixel = 59;
			6125: Pixel = 80;
			6126: Pixel = 140;
			6127: Pixel = 167;
			6128: Pixel = 176;
			6129: Pixel = 180;
			6130: Pixel = 180;
			6131: Pixel = 162;
			6132: Pixel = 121;
			6133: Pixel = 80;
			6134: Pixel = 86;
			6135: Pixel = 107;
			6136: Pixel = 124;
			6137: Pixel = 134;
			6138: Pixel = 123;
			6139: Pixel = 89;
			6140: Pixel = 74;
			6141: Pixel = 57;
			6142: Pixel = 66;
			6143: Pixel = 83;
			6144: Pixel = 103;
			6145: Pixel = 116;
			6146: Pixel = 79;
			6147: Pixel = 44;
			6148: Pixel = 46;
			6149: Pixel = 44;
			6150: Pixel = 67;
			6151: Pixel = 90;
			6152: Pixel = 55;
			6153: Pixel = 68;
			6154: Pixel = 135;
			6155: Pixel = 60;
			6156: Pixel = 43;
			6157: Pixel = 46;
			6158: Pixel = 41;
			6159: Pixel = 112;
			6160: Pixel = 141;
			6161: Pixel = 196;
			6162: Pixel = 172;
			6163: Pixel = 45;
			6164: Pixel = 88;
			6165: Pixel = 121;
			6166: Pixel = 125;
			6167: Pixel = 137;
			6168: Pixel = 148;
			6169: Pixel = 158;
			6170: Pixel = 171;
			6171: Pixel = 176;
			6172: Pixel = 178;
			6173: Pixel = 176;
			6174: Pixel = 175;
			6175: Pixel = 170;
			6176: Pixel = 156;
			6177: Pixel = 148;
			6178: Pixel = 141;
			6179: Pixel = 131;
			6180: Pixel = 128;
			6181: Pixel = 173;
			6182: Pixel = 222;
			6183: Pixel = 185;
			6184: Pixel = 161;
			6185: Pixel = 151;
			6186: Pixel = 135;
			6187: Pixel = 129;
			6188: Pixel = 121;
			6189: Pixel = 70;
			6190: Pixel = 50;
			6191: Pixel = 68;
			6192: Pixel = 47;
			6193: Pixel = 133;
			6194: Pixel = 143;
			6195: Pixel = 44;
			6196: Pixel = 49;
			6197: Pixel = 45;
			6198: Pixel = 67;
			6199: Pixel = 138;
			6200: Pixel = 142;
			6201: Pixel = 159;
			6202: Pixel = 154;
			6203: Pixel = 154;
			6204: Pixel = 151;
			6205: Pixel = 150;
			6206: Pixel = 150;
			6207: Pixel = 149;
			6208: Pixel = 147;
			6209: Pixel = 145;
			6210: Pixel = 145;
			6211: Pixel = 141;
			6212: Pixel = 133;
			6213: Pixel = 133;
			6214: Pixel = 174;
			6215: Pixel = 195;
			6216: Pixel = 194;
			6217: Pixel = 195;
			6218: Pixel = 193;
			6219: Pixel = 191;
			6220: Pixel = 194;
			6221: Pixel = 199;
			6222: Pixel = 79;
			6223: Pixel = 76;
			6224: Pixel = 74;
			6225: Pixel = 71;
			6226: Pixel = 58;
			6227: Pixel = 77;
			6228: Pixel = 139;
			6229: Pixel = 165;
			6230: Pixel = 175;
			6231: Pixel = 177;
			6232: Pixel = 177;
			6233: Pixel = 162;
			6234: Pixel = 122;
			6235: Pixel = 80;
			6236: Pixel = 88;
			6237: Pixel = 102;
			6238: Pixel = 106;
			6239: Pixel = 110;
			6240: Pixel = 98;
			6241: Pixel = 99;
			6242: Pixel = 90;
			6243: Pixel = 81;
			6244: Pixel = 90;
			6245: Pixel = 61;
			6246: Pixel = 108;
			6247: Pixel = 92;
			6248: Pixel = 56;
			6249: Pixel = 47;
			6250: Pixel = 51;
			6251: Pixel = 49;
			6252: Pixel = 50;
			6253: Pixel = 58;
			6254: Pixel = 43;
			6255: Pixel = 68;
			6256: Pixel = 134;
			6257: Pixel = 95;
			6258: Pixel = 32;
			6259: Pixel = 33;
			6260: Pixel = 69;
			6261: Pixel = 126;
			6262: Pixel = 172;
			6263: Pixel = 203;
			6264: Pixel = 74;
			6265: Pixel = 43;
			6266: Pixel = 97;
			6267: Pixel = 122;
			6268: Pixel = 127;
			6269: Pixel = 135;
			6270: Pixel = 145;
			6271: Pixel = 152;
			6272: Pixel = 163;
			6273: Pixel = 174;
			6274: Pixel = 179;
			6275: Pixel = 176;
			6276: Pixel = 171;
			6277: Pixel = 165;
			6278: Pixel = 151;
			6279: Pixel = 144;
			6280: Pixel = 141;
			6281: Pixel = 128;
			6282: Pixel = 130;
			6283: Pixel = 165;
			6284: Pixel = 220;
			6285: Pixel = 188;
			6286: Pixel = 159;
			6287: Pixel = 153;
			6288: Pixel = 139;
			6289: Pixel = 131;
			6290: Pixel = 117;
			6291: Pixel = 63;
			6292: Pixel = 46;
			6293: Pixel = 68;
			6294: Pixel = 43;
			6295: Pixel = 124;
			6296: Pixel = 155;
			6297: Pixel = 49;
			6298: Pixel = 51;
			6299: Pixel = 46;
			6300: Pixel = 89;
			6301: Pixel = 141;
			6302: Pixel = 153;
			6303: Pixel = 161;
			6304: Pixel = 153;
			6305: Pixel = 154;
			6306: Pixel = 151;
			6307: Pixel = 149;
			6308: Pixel = 147;
			6309: Pixel = 147;
			6310: Pixel = 146;
			6311: Pixel = 144;
			6312: Pixel = 143;
			6313: Pixel = 138;
			6314: Pixel = 128;
			6315: Pixel = 156;
			6316: Pixel = 194;
			6317: Pixel = 194;
			6318: Pixel = 192;
			6319: Pixel = 194;
			6320: Pixel = 194;
			6321: Pixel = 198;
			6322: Pixel = 203;
			6323: Pixel = 204;
			6324: Pixel = 76;
			6325: Pixel = 75;
			6326: Pixel = 74;
			6327: Pixel = 69;
			6328: Pixel = 53;
			6329: Pixel = 76;
			6330: Pixel = 139;
			6331: Pixel = 164;
			6332: Pixel = 173;
			6333: Pixel = 173;
			6334: Pixel = 175;
			6335: Pixel = 160;
			6336: Pixel = 123;
			6337: Pixel = 74;
			6338: Pixel = 100;
			6339: Pixel = 102;
			6340: Pixel = 116;
			6341: Pixel = 133;
			6342: Pixel = 98;
			6343: Pixel = 93;
			6344: Pixel = 110;
			6345: Pixel = 88;
			6346: Pixel = 69;
			6347: Pixel = 65;
			6348: Pixel = 100;
			6349: Pixel = 111;
			6350: Pixel = 59;
			6351: Pixel = 58;
			6352: Pixel = 50;
			6353: Pixel = 41;
			6354: Pixel = 50;
			6355: Pixel = 69;
			6356: Pixel = 46;
			6357: Pixel = 90;
			6358: Pixel = 115;
			6359: Pixel = 130;
			6360: Pixel = 70;
			6361: Pixel = 28;
			6362: Pixel = 103;
			6363: Pixel = 135;
			6364: Pixel = 214;
			6365: Pixel = 133;
			6366: Pixel = 32;
			6367: Pixel = 61;
			6368: Pixel = 89;
			6369: Pixel = 119;
			6370: Pixel = 128;
			6371: Pixel = 134;
			6372: Pixel = 144;
			6373: Pixel = 152;
			6374: Pixel = 157;
			6375: Pixel = 167;
			6376: Pixel = 174;
			6377: Pixel = 173;
			6378: Pixel = 169;
			6379: Pixel = 162;
			6380: Pixel = 147;
			6381: Pixel = 135;
			6382: Pixel = 134;
			6383: Pixel = 124;
			6384: Pixel = 128;
			6385: Pixel = 156;
			6386: Pixel = 215;
			6387: Pixel = 193;
			6388: Pixel = 155;
			6389: Pixel = 150;
			6390: Pixel = 139;
			6391: Pixel = 132;
			6392: Pixel = 109;
			6393: Pixel = 52;
			6394: Pixel = 49;
			6395: Pixel = 72;
			6396: Pixel = 39;
			6397: Pixel = 112;
			6398: Pixel = 160;
			6399: Pixel = 66;
			6400: Pixel = 46;
			6401: Pixel = 49;
			6402: Pixel = 113;
			6403: Pixel = 142;
			6404: Pixel = 159;
			6405: Pixel = 159;
			6406: Pixel = 154;
			6407: Pixel = 153;
			6408: Pixel = 151;
			6409: Pixel = 148;
			6410: Pixel = 146;
			6411: Pixel = 145;
			6412: Pixel = 143;
			6413: Pixel = 143;
			6414: Pixel = 141;
			6415: Pixel = 132;
			6416: Pixel = 138;
			6417: Pixel = 184;
			6418: Pixel = 196;
			6419: Pixel = 192;
			6420: Pixel = 192;
			6421: Pixel = 195;
			6422: Pixel = 202;
			6423: Pixel = 208;
			6424: Pixel = 205;
			6425: Pixel = 201;
			6426: Pixel = 78;
			6427: Pixel = 76;
			6428: Pixel = 74;
			6429: Pixel = 67;
			6430: Pixel = 50;
			6431: Pixel = 74;
			6432: Pixel = 138;
			6433: Pixel = 164;
			6434: Pixel = 172;
			6435: Pixel = 173;
			6436: Pixel = 175;
			6437: Pixel = 160;
			6438: Pixel = 121;
			6439: Pixel = 72;
			6440: Pixel = 95;
			6441: Pixel = 125;
			6442: Pixel = 131;
			6443: Pixel = 125;
			6444: Pixel = 63;
			6445: Pixel = 108;
			6446: Pixel = 100;
			6447: Pixel = 66;
			6448: Pixel = 82;
			6449: Pixel = 97;
			6450: Pixel = 114;
			6451: Pixel = 119;
			6452: Pixel = 72;
			6453: Pixel = 53;
			6454: Pixel = 46;
			6455: Pixel = 36;
			6456: Pixel = 63;
			6457: Pixel = 91;
			6458: Pixel = 67;
			6459: Pixel = 126;
			6460: Pixel = 152;
			6461: Pixel = 76;
			6462: Pixel = 56;
			6463: Pixel = 47;
			6464: Pixel = 124;
			6465: Pixel = 175;
			6466: Pixel = 183;
			6467: Pixel = 38;
			6468: Pixel = 44;
			6469: Pixel = 67;
			6470: Pixel = 85;
			6471: Pixel = 117;
			6472: Pixel = 127;
			6473: Pixel = 132;
			6474: Pixel = 140;
			6475: Pixel = 149;
			6476: Pixel = 156;
			6477: Pixel = 159;
			6478: Pixel = 164;
			6479: Pixel = 167;
			6480: Pixel = 166;
			6481: Pixel = 160;
			6482: Pixel = 144;
			6483: Pixel = 131;
			6484: Pixel = 129;
			6485: Pixel = 122;
			6486: Pixel = 123;
			6487: Pixel = 149;
			6488: Pixel = 208;
			6489: Pixel = 204;
			6490: Pixel = 153;
			6491: Pixel = 149;
			6492: Pixel = 137;
			6493: Pixel = 131;
			6494: Pixel = 94;
			6495: Pixel = 43;
			6496: Pixel = 55;
			6497: Pixel = 76;
			6498: Pixel = 39;
			6499: Pixel = 99;
			6500: Pixel = 164;
			6501: Pixel = 75;
			6502: Pixel = 37;
			6503: Pixel = 58;
			6504: Pixel = 131;
			6505: Pixel = 144;
			6506: Pixel = 159;
			6507: Pixel = 156;
			6508: Pixel = 152;
			6509: Pixel = 154;
			6510: Pixel = 152;
			6511: Pixel = 149;
			6512: Pixel = 147;
			6513: Pixel = 146;
			6514: Pixel = 144;
			6515: Pixel = 141;
			6516: Pixel = 138;
			6517: Pixel = 130;
			6518: Pixel = 162;
			6519: Pixel = 196;
			6520: Pixel = 194;
			6521: Pixel = 192;
			6522: Pixel = 194;
			6523: Pixel = 204;
			6524: Pixel = 207;
			6525: Pixel = 209;
			6526: Pixel = 205;
			6527: Pixel = 203;
			6528: Pixel = 80;
			6529: Pixel = 76;
			6530: Pixel = 74;
			6531: Pixel = 64;
			6532: Pixel = 45;
			6533: Pixel = 67;
			6534: Pixel = 136;
			6535: Pixel = 164;
			6536: Pixel = 173;
			6537: Pixel = 175;
			6538: Pixel = 177;
			6539: Pixel = 162;
			6540: Pixel = 122;
			6541: Pixel = 73;
			6542: Pixel = 84;
			6543: Pixel = 116;
			6544: Pixel = 116;
			6545: Pixel = 114;
			6546: Pixel = 75;
			6547: Pixel = 92;
			6548: Pixel = 90;
			6549: Pixel = 76;
			6550: Pixel = 92;
			6551: Pixel = 85;
			6552: Pixel = 103;
			6553: Pixel = 118;
			6554: Pixel = 64;
			6555: Pixel = 42;
			6556: Pixel = 54;
			6557: Pixel = 41;
			6558: Pixel = 66;
			6559: Pixel = 87;
			6560: Pixel = 123;
			6561: Pixel = 97;
			6562: Pixel = 87;
			6563: Pixel = 42;
			6564: Pixel = 38;
			6565: Pixel = 96;
			6566: Pixel = 124;
			6567: Pixel = 189;
			6568: Pixel = 83;
			6569: Pixel = 24;
			6570: Pixel = 54;
			6571: Pixel = 78;
			6572: Pixel = 83;
			6573: Pixel = 115;
			6574: Pixel = 125;
			6575: Pixel = 132;
			6576: Pixel = 137;
			6577: Pixel = 145;
			6578: Pixel = 151;
			6579: Pixel = 153;
			6580: Pixel = 157;
			6581: Pixel = 162;
			6582: Pixel = 161;
			6583: Pixel = 154;
			6584: Pixel = 136;
			6585: Pixel = 120;
			6586: Pixel = 134;
			6587: Pixel = 130;
			6588: Pixel = 124;
			6589: Pixel = 144;
			6590: Pixel = 200;
			6591: Pixel = 214;
			6592: Pixel = 149;
			6593: Pixel = 149;
			6594: Pixel = 135;
			6595: Pixel = 128;
			6596: Pixel = 74;
			6597: Pixel = 40;
			6598: Pixel = 58;
			6599: Pixel = 75;
			6600: Pixel = 38;
			6601: Pixel = 84;
			6602: Pixel = 167;
			6603: Pixel = 96;
			6604: Pixel = 30;
			6605: Pixel = 80;
			6606: Pixel = 142;
			6607: Pixel = 147;
			6608: Pixel = 159;
			6609: Pixel = 154;
			6610: Pixel = 151;
			6611: Pixel = 150;
			6612: Pixel = 151;
			6613: Pixel = 150;
			6614: Pixel = 148;
			6615: Pixel = 147;
			6616: Pixel = 145;
			6617: Pixel = 142;
			6618: Pixel = 133;
			6619: Pixel = 139;
			6620: Pixel = 187;
			6621: Pixel = 197;
			6622: Pixel = 193;
			6623: Pixel = 194;
			6624: Pixel = 203;
			6625: Pixel = 208;
			6626: Pixel = 205;
			6627: Pixel = 205;
			6628: Pixel = 207;
			6629: Pixel = 207;
			6630: Pixel = 84;
			6631: Pixel = 80;
			6632: Pixel = 74;
			6633: Pixel = 66;
			6634: Pixel = 46;
			6635: Pixel = 69;
			6636: Pixel = 136;
			6637: Pixel = 165;
			6638: Pixel = 173;
			6639: Pixel = 175;
			6640: Pixel = 178;
			6641: Pixel = 163;
			6642: Pixel = 122;
			6643: Pixel = 86;
			6644: Pixel = 111;
			6645: Pixel = 107;
			6646: Pixel = 114;
			6647: Pixel = 99;
			6648: Pixel = 68;
			6649: Pixel = 104;
			6650: Pixel = 91;
			6651: Pixel = 64;
			6652: Pixel = 94;
			6653: Pixel = 65;
			6654: Pixel = 102;
			6655: Pixel = 116;
			6656: Pixel = 81;
			6657: Pixel = 59;
			6658: Pixel = 56;
			6659: Pixel = 43;
			6660: Pixel = 60;
			6661: Pixel = 80;
			6662: Pixel = 82;
			6663: Pixel = 90;
			6664: Pixel = 37;
			6665: Pixel = 26;
			6666: Pixel = 105;
			6667: Pixel = 167;
			6668: Pixel = 154;
			6669: Pixel = 148;
			6670: Pixel = 45;
			6671: Pixel = 37;
			6672: Pixel = 56;
			6673: Pixel = 85;
			6674: Pixel = 83;
			6675: Pixel = 116;
			6676: Pixel = 126;
			6677: Pixel = 129;
			6678: Pixel = 138;
			6679: Pixel = 143;
			6680: Pixel = 148;
			6681: Pixel = 152;
			6682: Pixel = 155;
			6683: Pixel = 158;
			6684: Pixel = 159;
			6685: Pixel = 152;
			6686: Pixel = 130;
			6687: Pixel = 121;
			6688: Pixel = 134;
			6689: Pixel = 131;
			6690: Pixel = 126;
			6691: Pixel = 136;
			6692: Pixel = 194;
			6693: Pixel = 202;
			6694: Pixel = 145;
			6695: Pixel = 144;
			6696: Pixel = 134;
			6697: Pixel = 114;
			6698: Pixel = 49;
			6699: Pixel = 43;
			6700: Pixel = 59;
			6701: Pixel = 72;
			6702: Pixel = 41;
			6703: Pixel = 68;
			6704: Pixel = 167;
			6705: Pixel = 113;
			6706: Pixel = 29;
			6707: Pixel = 99;
			6708: Pixel = 149;
			6709: Pixel = 151;
			6710: Pixel = 157;
			6711: Pixel = 153;
			6712: Pixel = 150;
			6713: Pixel = 150;
			6714: Pixel = 149;
			6715: Pixel = 149;
			6716: Pixel = 148;
			6717: Pixel = 147;
			6718: Pixel = 145;
			6719: Pixel = 140;
			6720: Pixel = 129;
			6721: Pixel = 158;
			6722: Pixel = 196;
			6723: Pixel = 194;
			6724: Pixel = 193;
			6725: Pixel = 199;
			6726: Pixel = 206;
			6727: Pixel = 206;
			6728: Pixel = 204;
			6729: Pixel = 205;
			6730: Pixel = 208;
			6731: Pixel = 207;
			6732: Pixel = 81;
			6733: Pixel = 78;
			6734: Pixel = 76;
			6735: Pixel = 69;
			6736: Pixel = 56;
			6737: Pixel = 85;
			6738: Pixel = 142;
			6739: Pixel = 164;
			6740: Pixel = 172;
			6741: Pixel = 175;
			6742: Pixel = 178;
			6743: Pixel = 163;
			6744: Pixel = 127;
			6745: Pixel = 85;
			6746: Pixel = 84;
			6747: Pixel = 96;
			6748: Pixel = 113;
			6749: Pixel = 94;
			6750: Pixel = 77;
			6751: Pixel = 112;
			6752: Pixel = 72;
			6753: Pixel = 75;
			6754: Pixel = 101;
			6755: Pixel = 65;
			6756: Pixel = 96;
			6757: Pixel = 128;
			6758: Pixel = 103;
			6759: Pixel = 58;
			6760: Pixel = 57;
			6761: Pixel = 61;
			6762: Pixel = 35;
			6763: Pixel = 48;
			6764: Pixel = 104;
			6765: Pixel = 55;
			6766: Pixel = 37;
			6767: Pixel = 36;
			6768: Pixel = 147;
			6769: Pixel = 191;
			6770: Pixel = 177;
			6771: Pixel = 56;
			6772: Pixel = 35;
			6773: Pixel = 43;
			6774: Pixel = 55;
			6775: Pixel = 92;
			6776: Pixel = 91;
			6777: Pixel = 115;
			6778: Pixel = 124;
			6779: Pixel = 129;
			6780: Pixel = 136;
			6781: Pixel = 143;
			6782: Pixel = 148;
			6783: Pixel = 150;
			6784: Pixel = 152;
			6785: Pixel = 156;
			6786: Pixel = 158;
			6787: Pixel = 154;
			6788: Pixel = 138;
			6789: Pixel = 128;
			6790: Pixel = 107;
			6791: Pixel = 90;
			6792: Pixel = 107;
			6793: Pixel = 113;
			6794: Pixel = 168;
			6795: Pixel = 177;
			6796: Pixel = 146;
			6797: Pixel = 141;
			6798: Pixel = 135;
			6799: Pixel = 85;
			6800: Pixel = 40;
			6801: Pixel = 49;
			6802: Pixel = 62;
			6803: Pixel = 68;
			6804: Pixel = 47;
			6805: Pixel = 55;
			6806: Pixel = 158;
			6807: Pixel = 119;
			6808: Pixel = 45;
			6809: Pixel = 122;
			6810: Pixel = 149;
			6811: Pixel = 154;
			6812: Pixel = 155;
			6813: Pixel = 151;
			6814: Pixel = 150;
			6815: Pixel = 150;
			6816: Pixel = 150;
			6817: Pixel = 147;
			6818: Pixel = 146;
			6819: Pixel = 144;
			6820: Pixel = 144;
			6821: Pixel = 138;
			6822: Pixel = 133;
			6823: Pixel = 174;
			6824: Pixel = 198;
			6825: Pixel = 194;
			6826: Pixel = 198;
			6827: Pixel = 206;
			6828: Pixel = 205;
			6829: Pixel = 206;
			6830: Pixel = 209;
			6831: Pixel = 209;
			6832: Pixel = 209;
			6833: Pixel = 206;
			6834: Pixel = 79;
			6835: Pixel = 77;
			6836: Pixel = 75;
			6837: Pixel = 69;
			6838: Pixel = 70;
			6839: Pixel = 103;
			6840: Pixel = 149;
			6841: Pixel = 164;
			6842: Pixel = 170;
			6843: Pixel = 173;
			6844: Pixel = 179;
			6845: Pixel = 165;
			6846: Pixel = 126;
			6847: Pixel = 77;
			6848: Pixel = 85;
			6849: Pixel = 99;
			6850: Pixel = 116;
			6851: Pixel = 87;
			6852: Pixel = 70;
			6853: Pixel = 75;
			6854: Pixel = 60;
			6855: Pixel = 96;
			6856: Pixel = 77;
			6857: Pixel = 81;
			6858: Pixel = 98;
			6859: Pixel = 114;
			6860: Pixel = 130;
			6861: Pixel = 68;
			6862: Pixel = 37;
			6863: Pixel = 128;
			6864: Pixel = 55;
			6865: Pixel = 53;
			6866: Pixel = 81;
			6867: Pixel = 58;
			6868: Pixel = 100;
			6869: Pixel = 120;
			6870: Pixel = 113;
			6871: Pixel = 174;
			6872: Pixel = 86;
			6873: Pixel = 32;
			6874: Pixel = 62;
			6875: Pixel = 42;
			6876: Pixel = 59;
			6877: Pixel = 100;
			6878: Pixel = 95;
			6879: Pixel = 118;
			6880: Pixel = 123;
			6881: Pixel = 128;
			6882: Pixel = 133;
			6883: Pixel = 141;
			6884: Pixel = 146;
			6885: Pixel = 146;
			6886: Pixel = 151;
			6887: Pixel = 154;
			6888: Pixel = 158;
			6889: Pixel = 156;
			6890: Pixel = 150;
			6891: Pixel = 136;
			6892: Pixel = 129;
			6893: Pixel = 135;
			6894: Pixel = 126;
			6895: Pixel = 151;
			6896: Pixel = 183;
			6897: Pixel = 167;
			6898: Pixel = 148;
			6899: Pixel = 138;
			6900: Pixel = 124;
			6901: Pixel = 56;
			6902: Pixel = 46;
			6903: Pixel = 50;
			6904: Pixel = 70;
			6905: Pixel = 74;
			6906: Pixel = 52;
			6907: Pixel = 45;
			6908: Pixel = 146;
			6909: Pixel = 125;
			6910: Pixel = 64;
			6911: Pixel = 139;
			6912: Pixel = 149;
			6913: Pixel = 156;
			6914: Pixel = 154;
			6915: Pixel = 151;
			6916: Pixel = 150;
			6917: Pixel = 149;
			6918: Pixel = 149;
			6919: Pixel = 148;
			6920: Pixel = 145;
			6921: Pixel = 144;
			6922: Pixel = 143;
			6923: Pixel = 135;
			6924: Pixel = 140;
			6925: Pixel = 185;
			6926: Pixel = 196;
			6927: Pixel = 196;
			6928: Pixel = 204;
			6929: Pixel = 207;
			6930: Pixel = 206;
			6931: Pixel = 207;
			6932: Pixel = 210;
			6933: Pixel = 209;
			6934: Pixel = 207;
			6935: Pixel = 207;
			6936: Pixel = 77;
			6937: Pixel = 76;
			6938: Pixel = 78;
			6939: Pixel = 67;
			6940: Pixel = 70;
			6941: Pixel = 113;
			6942: Pixel = 152;
			6943: Pixel = 164;
			6944: Pixel = 169;
			6945: Pixel = 174;
			6946: Pixel = 179;
			6947: Pixel = 165;
			6948: Pixel = 128;
			6949: Pixel = 80;
			6950: Pixel = 85;
			6951: Pixel = 94;
			6952: Pixel = 129;
			6953: Pixel = 98;
			6954: Pixel = 55;
			6955: Pixel = 82;
			6956: Pixel = 100;
			6957: Pixel = 56;
			6958: Pixel = 63;
			6959: Pixel = 83;
			6960: Pixel = 104;
			6961: Pixel = 100;
			6962: Pixel = 125;
			6963: Pixel = 109;
			6964: Pixel = 54;
			6965: Pixel = 107;
			6966: Pixel = 73;
			6967: Pixel = 44;
			6968: Pixel = 86;
			6969: Pixel = 132;
			6970: Pixel = 170;
			6971: Pixel = 115;
			6972: Pixel = 130;
			6973: Pixel = 138;
			6974: Pixel = 38;
			6975: Pixel = 54;
			6976: Pixel = 59;
			6977: Pixel = 50;
			6978: Pixel = 58;
			6979: Pixel = 103;
			6980: Pixel = 98;
			6981: Pixel = 120;
			6982: Pixel = 125;
			6983: Pixel = 127;
			6984: Pixel = 134;
			6985: Pixel = 140;
			6986: Pixel = 142;
			6987: Pixel = 144;
			6988: Pixel = 151;
			6989: Pixel = 154;
			6990: Pixel = 157;
			6991: Pixel = 156;
			6992: Pixel = 152;
			6993: Pixel = 149;
			6994: Pixel = 141;
			6995: Pixel = 162;
			6996: Pixel = 176;
			6997: Pixel = 189;
			6998: Pixel = 196;
			6999: Pixel = 162;
			7000: Pixel = 144;
			7001: Pixel = 141;
			7002: Pixel = 96;
			7003: Pixel = 45;
			7004: Pixel = 47;
			7005: Pixel = 56;
			7006: Pixel = 76;
			7007: Pixel = 74;
			7008: Pixel = 61;
			7009: Pixel = 40;
			7010: Pixel = 132;
			7011: Pixel = 127;
			7012: Pixel = 91;
			7013: Pixel = 145;
			7014: Pixel = 149;
			7015: Pixel = 156;
			7016: Pixel = 153;
			7017: Pixel = 151;
			7018: Pixel = 150;
			7019: Pixel = 148;
			7020: Pixel = 147;
			7021: Pixel = 146;
			7022: Pixel = 146;
			7023: Pixel = 144;
			7024: Pixel = 142;
			7025: Pixel = 132;
			7026: Pixel = 147;
			7027: Pixel = 191;
			7028: Pixel = 195;
			7029: Pixel = 200;
			7030: Pixel = 208;
			7031: Pixel = 207;
			7032: Pixel = 205;
			7033: Pixel = 208;
			7034: Pixel = 208;
			7035: Pixel = 210;
			7036: Pixel = 210;
			7037: Pixel = 210;
			7038: Pixel = 73;
			7039: Pixel = 71;
			7040: Pixel = 72;
			7041: Pixel = 64;
			7042: Pixel = 69;
			7043: Pixel = 114;
			7044: Pixel = 151;
			7045: Pixel = 165;
			7046: Pixel = 169;
			7047: Pixel = 174;
			7048: Pixel = 179;
			7049: Pixel = 166;
			7050: Pixel = 128;
			7051: Pixel = 79;
			7052: Pixel = 78;
			7053: Pixel = 107;
			7054: Pixel = 134;
			7055: Pixel = 87;
			7056: Pixel = 75;
			7057: Pixel = 108;
			7058: Pixel = 62;
			7059: Pixel = 58;
			7060: Pixel = 64;
			7061: Pixel = 69;
			7062: Pixel = 81;
			7063: Pixel = 88;
			7064: Pixel = 105;
			7065: Pixel = 126;
			7066: Pixel = 99;
			7067: Pixel = 79;
			7068: Pixel = 46;
			7069: Pixel = 63;
			7070: Pixel = 126;
			7071: Pixel = 180;
			7072: Pixel = 156;
			7073: Pixel = 87;
			7074: Pixel = 136;
			7075: Pixel = 47;
			7076: Pixel = 47;
			7077: Pixel = 48;
			7078: Pixel = 60;
			7079: Pixel = 55;
			7080: Pixel = 50;
			7081: Pixel = 101;
			7082: Pixel = 100;
			7083: Pixel = 117;
			7084: Pixel = 126;
			7085: Pixel = 128;
			7086: Pixel = 134;
			7087: Pixel = 140;
			7088: Pixel = 140;
			7089: Pixel = 140;
			7090: Pixel = 144;
			7091: Pixel = 149;
			7092: Pixel = 149;
			7093: Pixel = 152;
			7094: Pixel = 148;
			7095: Pixel = 149;
			7096: Pixel = 149;
			7097: Pixel = 186;
			7098: Pixel = 197;
			7099: Pixel = 188;
			7100: Pixel = 199;
			7101: Pixel = 158;
			7102: Pixel = 142;
			7103: Pixel = 135;
			7104: Pixel = 61;
			7105: Pixel = 45;
			7106: Pixel = 48;
			7107: Pixel = 60;
			7108: Pixel = 76;
			7109: Pixel = 70;
			7110: Pixel = 60;
			7111: Pixel = 36;
			7112: Pixel = 118;
			7113: Pixel = 130;
			7114: Pixel = 113;
			7115: Pixel = 147;
			7116: Pixel = 151;
			7117: Pixel = 155;
			7118: Pixel = 152;
			7119: Pixel = 150;
			7120: Pixel = 148;
			7121: Pixel = 148;
			7122: Pixel = 146;
			7123: Pixel = 144;
			7124: Pixel = 145;
			7125: Pixel = 144;
			7126: Pixel = 141;
			7127: Pixel = 130;
			7128: Pixel = 154;
			7129: Pixel = 194;
			7130: Pixel = 197;
			7131: Pixel = 206;
			7132: Pixel = 209;
			7133: Pixel = 206;
			7134: Pixel = 207;
			7135: Pixel = 207;
			7136: Pixel = 208;
			7137: Pixel = 211;
			7138: Pixel = 210;
			7139: Pixel = 211;
			7140: Pixel = 68;
			7141: Pixel = 66;
			7142: Pixel = 69;
			7143: Pixel = 64;
			7144: Pixel = 70;
			7145: Pixel = 108;
			7146: Pixel = 150;
			7147: Pixel = 165;
			7148: Pixel = 170;
			7149: Pixel = 175;
			7150: Pixel = 180;
			7151: Pixel = 168;
			7152: Pixel = 129;
			7153: Pixel = 75;
			7154: Pixel = 85;
			7155: Pixel = 120;
			7156: Pixel = 112;
			7157: Pixel = 84;
			7158: Pixel = 82;
			7159: Pixel = 89;
			7160: Pixel = 50;
			7161: Pixel = 70;
			7162: Pixel = 71;
			7163: Pixel = 80;
			7164: Pixel = 71;
			7165: Pixel = 81;
			7166: Pixel = 76;
			7167: Pixel = 117;
			7168: Pixel = 129;
			7169: Pixel = 40;
			7170: Pixel = 89;
			7171: Pixel = 136;
			7172: Pixel = 151;
			7173: Pixel = 178;
			7174: Pixel = 95;
			7175: Pixel = 130;
			7176: Pixel = 67;
			7177: Pixel = 51;
			7178: Pixel = 62;
			7179: Pixel = 46;
			7180: Pixel = 62;
			7181: Pixel = 62;
			7182: Pixel = 45;
			7183: Pixel = 95;
			7184: Pixel = 93;
			7185: Pixel = 112;
			7186: Pixel = 126;
			7187: Pixel = 128;
			7188: Pixel = 133;
			7189: Pixel = 139;
			7190: Pixel = 140;
			7191: Pixel = 137;
			7192: Pixel = 140;
			7193: Pixel = 144;
			7194: Pixel = 145;
			7195: Pixel = 146;
			7196: Pixel = 146;
			7197: Pixel = 151;
			7198: Pixel = 158;
			7199: Pixel = 175;
			7200: Pixel = 192;
			7201: Pixel = 190;
			7202: Pixel = 186;
			7203: Pixel = 147;
			7204: Pixel = 140;
			7205: Pixel = 109;
			7206: Pixel = 41;
			7207: Pixel = 53;
			7208: Pixel = 49;
			7209: Pixel = 61;
			7210: Pixel = 77;
			7211: Pixel = 71;
			7212: Pixel = 63;
			7213: Pixel = 34;
			7214: Pixel = 108;
			7215: Pixel = 135;
			7216: Pixel = 123;
			7217: Pixel = 146;
			7218: Pixel = 152;
			7219: Pixel = 154;
			7220: Pixel = 152;
			7221: Pixel = 150;
			7222: Pixel = 147;
			7223: Pixel = 148;
			7224: Pixel = 147;
			7225: Pixel = 145;
			7226: Pixel = 145;
			7227: Pixel = 143;
			7228: Pixel = 139;
			7229: Pixel = 128;
			7230: Pixel = 158;
			7231: Pixel = 196;
			7232: Pixel = 202;
			7233: Pixel = 209;
			7234: Pixel = 207;
			7235: Pixel = 208;
			7236: Pixel = 208;
			7237: Pixel = 207;
			7238: Pixel = 211;
			7239: Pixel = 212;
			7240: Pixel = 211;
			7241: Pixel = 211;
			7242: Pixel = 59;
			7243: Pixel = 59;
			7244: Pixel = 66;
			7245: Pixel = 63;
			7246: Pixel = 69;
			7247: Pixel = 109;
			7248: Pixel = 152;
			7249: Pixel = 167;
			7250: Pixel = 173;
			7251: Pixel = 176;
			7252: Pixel = 180;
			7253: Pixel = 168;
			7254: Pixel = 126;
			7255: Pixel = 72;
			7256: Pixel = 113;
			7257: Pixel = 97;
			7258: Pixel = 125;
			7259: Pixel = 77;
			7260: Pixel = 61;
			7261: Pixel = 75;
			7262: Pixel = 64;
			7263: Pixel = 59;
			7264: Pixel = 68;
			7265: Pixel = 108;
			7266: Pixel = 95;
			7267: Pixel = 77;
			7268: Pixel = 83;
			7269: Pixel = 93;
			7270: Pixel = 103;
			7271: Pixel = 92;
			7272: Pixel = 131;
			7273: Pixel = 189;
			7274: Pixel = 207;
			7275: Pixel = 109;
			7276: Pixel = 116;
			7277: Pixel = 111;
			7278: Pixel = 30;
			7279: Pixel = 61;
			7280: Pixel = 57;
			7281: Pixel = 44;
			7282: Pixel = 63;
			7283: Pixel = 66;
			7284: Pixel = 46;
			7285: Pixel = 89;
			7286: Pixel = 84;
			7287: Pixel = 104;
			7288: Pixel = 126;
			7289: Pixel = 129;
			7290: Pixel = 129;
			7291: Pixel = 135;
			7292: Pixel = 140;
			7293: Pixel = 142;
			7294: Pixel = 135;
			7295: Pixel = 105;
			7296: Pixel = 112;
			7297: Pixel = 124;
			7298: Pixel = 126;
			7299: Pixel = 120;
			7300: Pixel = 112;
			7301: Pixel = 111;
			7302: Pixel = 130;
			7303: Pixel = 118;
			7304: Pixel = 115;
			7305: Pixel = 118;
			7306: Pixel = 142;
			7307: Pixel = 68;
			7308: Pixel = 43;
			7309: Pixel = 51;
			7310: Pixel = 51;
			7311: Pixel = 65;
			7312: Pixel = 74;
			7313: Pixel = 74;
			7314: Pixel = 63;
			7315: Pixel = 37;
			7316: Pixel = 92;
			7317: Pixel = 140;
			7318: Pixel = 135;
			7319: Pixel = 147;
			7320: Pixel = 153;
			7321: Pixel = 155;
			7322: Pixel = 151;
			7323: Pixel = 149;
			7324: Pixel = 147;
			7325: Pixel = 148;
			7326: Pixel = 147;
			7327: Pixel = 145;
			7328: Pixel = 143;
			7329: Pixel = 143;
			7330: Pixel = 139;
			7331: Pixel = 127;
			7332: Pixel = 163;
			7333: Pixel = 200;
			7334: Pixel = 208;
			7335: Pixel = 210;
			7336: Pixel = 208;
			7337: Pixel = 208;
			7338: Pixel = 208;
			7339: Pixel = 210;
			7340: Pixel = 212;
			7341: Pixel = 213;
			7342: Pixel = 212;
			7343: Pixel = 212;
			7344: Pixel = 55;
			7345: Pixel = 59;
			7346: Pixel = 64;
			7347: Pixel = 62;
			7348: Pixel = 78;
			7349: Pixel = 115;
			7350: Pixel = 152;
			7351: Pixel = 169;
			7352: Pixel = 176;
			7353: Pixel = 178;
			7354: Pixel = 180;
			7355: Pixel = 165;
			7356: Pixel = 121;
			7357: Pixel = 115;
			7358: Pixel = 100;
			7359: Pixel = 99;
			7360: Pixel = 139;
			7361: Pixel = 75;
			7362: Pixel = 59;
			7363: Pixel = 49;
			7364: Pixel = 63;
			7365: Pixel = 65;
			7366: Pixel = 72;
			7367: Pixel = 125;
			7368: Pixel = 95;
			7369: Pixel = 100;
			7370: Pixel = 91;
			7371: Pixel = 99;
			7372: Pixel = 70;
			7373: Pixel = 121;
			7374: Pixel = 135;
			7375: Pixel = 199;
			7376: Pixel = 155;
			7377: Pixel = 98;
			7378: Pixel = 148;
			7379: Pixel = 51;
			7380: Pixel = 47;
			7381: Pixel = 48;
			7382: Pixel = 55;
			7383: Pixel = 49;
			7384: Pixel = 59;
			7385: Pixel = 66;
			7386: Pixel = 50;
			7387: Pixel = 80;
			7388: Pixel = 81;
			7389: Pixel = 98;
			7390: Pixel = 121;
			7391: Pixel = 125;
			7392: Pixel = 126;
			7393: Pixel = 132;
			7394: Pixel = 138;
			7395: Pixel = 147;
			7396: Pixel = 140;
			7397: Pixel = 118;
			7398: Pixel = 108;
			7399: Pixel = 108;
			7400: Pixel = 117;
			7401: Pixel = 122;
			7402: Pixel = 126;
			7403: Pixel = 135;
			7404: Pixel = 157;
			7405: Pixel = 137;
			7406: Pixel = 124;
			7407: Pixel = 145;
			7408: Pixel = 112;
			7409: Pixel = 41;
			7410: Pixel = 51;
			7411: Pixel = 47;
			7412: Pixel = 54;
			7413: Pixel = 63;
			7414: Pixel = 75;
			7415: Pixel = 71;
			7416: Pixel = 65;
			7417: Pixel = 50;
			7418: Pixel = 77;
			7419: Pixel = 150;
			7420: Pixel = 144;
			7421: Pixel = 149;
			7422: Pixel = 155;
			7423: Pixel = 153;
			7424: Pixel = 152;
			7425: Pixel = 152;
			7426: Pixel = 149;
			7427: Pixel = 146;
			7428: Pixel = 146;
			7429: Pixel = 146;
			7430: Pixel = 144;
			7431: Pixel = 144;
			7432: Pixel = 137;
			7433: Pixel = 127;
			7434: Pixel = 170;
			7435: Pixel = 206;
			7436: Pixel = 211;
			7437: Pixel = 210;
			7438: Pixel = 209;
			7439: Pixel = 208;
			7440: Pixel = 210;
			7441: Pixel = 211;
			7442: Pixel = 212;
			7443: Pixel = 213;
			7444: Pixel = 213;
			7445: Pixel = 212;
			7446: Pixel = 55;
			7447: Pixel = 57;
			7448: Pixel = 61;
			7449: Pixel = 59;
			7450: Pixel = 81;
			7451: Pixel = 113;
			7452: Pixel = 151;
			7453: Pixel = 167;
			7454: Pixel = 176;
			7455: Pixel = 179;
			7456: Pixel = 180;
			7457: Pixel = 167;
			7458: Pixel = 143;
			7459: Pixel = 102;
			7460: Pixel = 72;
			7461: Pixel = 127;
			7462: Pixel = 110;
			7463: Pixel = 75;
			7464: Pixel = 89;
			7465: Pixel = 46;
			7466: Pixel = 59;
			7467: Pixel = 75;
			7468: Pixel = 86;
			7469: Pixel = 133;
			7470: Pixel = 68;
			7471: Pixel = 97;
			7472: Pixel = 101;
			7473: Pixel = 73;
			7474: Pixel = 110;
			7475: Pixel = 147;
			7476: Pixel = 134;
			7477: Pixel = 163;
			7478: Pixel = 117;
			7479: Pixel = 162;
			7480: Pixel = 77;
			7481: Pixel = 45;
			7482: Pixel = 54;
			7483: Pixel = 45;
			7484: Pixel = 52;
			7485: Pixel = 49;
			7486: Pixel = 58;
			7487: Pixel = 65;
			7488: Pixel = 54;
			7489: Pixel = 73;
			7490: Pixel = 74;
			7491: Pixel = 88;
			7492: Pixel = 113;
			7493: Pixel = 118;
			7494: Pixel = 122;
			7495: Pixel = 126;
			7496: Pixel = 132;
			7497: Pixel = 141;
			7498: Pixel = 147;
			7499: Pixel = 141;
			7500: Pixel = 130;
			7501: Pixel = 127;
			7502: Pixel = 128;
			7503: Pixel = 139;
			7504: Pixel = 164;
			7505: Pixel = 170;
			7506: Pixel = 173;
			7507: Pixel = 151;
			7508: Pixel = 146;
			7509: Pixel = 143;
			7510: Pixel = 60;
			7511: Pixel = 43;
			7512: Pixel = 51;
			7513: Pixel = 44;
			7514: Pixel = 53;
			7515: Pixel = 58;
			7516: Pixel = 81;
			7517: Pixel = 73;
			7518: Pixel = 69;
			7519: Pixel = 54;
			7520: Pixel = 74;
			7521: Pixel = 156;
			7522: Pixel = 149;
			7523: Pixel = 150;
			7524: Pixel = 155;
			7525: Pixel = 154;
			7526: Pixel = 153;
			7527: Pixel = 152;
			7528: Pixel = 151;
			7529: Pixel = 149;
			7530: Pixel = 147;
			7531: Pixel = 145;
			7532: Pixel = 145;
			7533: Pixel = 144;
			7534: Pixel = 136;
			7535: Pixel = 126;
			7536: Pixel = 177;
			7537: Pixel = 213;
			7538: Pixel = 212;
			7539: Pixel = 210;
			7540: Pixel = 211;
			7541: Pixel = 211;
			7542: Pixel = 212;
			7543: Pixel = 214;
			7544: Pixel = 213;
			7545: Pixel = 209;
			7546: Pixel = 208;
			7547: Pixel = 207;
			7548: Pixel = 52;
			7549: Pixel = 53;
			7550: Pixel = 56;
			7551: Pixel = 56;
			7552: Pixel = 81;
			7553: Pixel = 106;
			7554: Pixel = 148;
			7555: Pixel = 165;
			7556: Pixel = 178;
			7557: Pixel = 179;
			7558: Pixel = 180;
			7559: Pixel = 169;
			7560: Pixel = 130;
			7561: Pixel = 63;
			7562: Pixel = 101;
			7563: Pixel = 125;
			7564: Pixel = 92;
			7565: Pixel = 71;
			7566: Pixel = 102;
			7567: Pixel = 39;
			7568: Pixel = 76;
			7569: Pixel = 65;
			7570: Pixel = 110;
			7571: Pixel = 125;
			7572: Pixel = 100;
			7573: Pixel = 85;
			7574: Pixel = 90;
			7575: Pixel = 124;
			7576: Pixel = 116;
			7577: Pixel = 140;
			7578: Pixel = 141;
			7579: Pixel = 159;
			7580: Pixel = 171;
			7581: Pixel = 105;
			7582: Pixel = 42;
			7583: Pixel = 57;
			7584: Pixel = 57;
			7585: Pixel = 51;
			7586: Pixel = 52;
			7587: Pixel = 55;
			7588: Pixel = 59;
			7589: Pixel = 66;
			7590: Pixel = 56;
			7591: Pixel = 72;
			7592: Pixel = 72;
			7593: Pixel = 75;
			7594: Pixel = 102;
			7595: Pixel = 109;
			7596: Pixel = 116;
			7597: Pixel = 124;
			7598: Pixel = 131;
			7599: Pixel = 135;
			7600: Pixel = 141;
			7601: Pixel = 141;
			7602: Pixel = 133;
			7603: Pixel = 128;
			7604: Pixel = 125;
			7605: Pixel = 121;
			7606: Pixel = 125;
			7607: Pixel = 127;
			7608: Pixel = 127;
			7609: Pixel = 142;
			7610: Pixel = 149;
			7611: Pixel = 99;
			7612: Pixel = 42;
			7613: Pixel = 46;
			7614: Pixel = 51;
			7615: Pixel = 54;
			7616: Pixel = 53;
			7617: Pixel = 61;
			7618: Pixel = 80;
			7619: Pixel = 76;
			7620: Pixel = 69;
			7621: Pixel = 59;
			7622: Pixel = 73;
			7623: Pixel = 158;
			7624: Pixel = 151;
			7625: Pixel = 151;
			7626: Pixel = 154;
			7627: Pixel = 153;
			7628: Pixel = 153;
			7629: Pixel = 153;
			7630: Pixel = 152;
			7631: Pixel = 150;
			7632: Pixel = 148;
			7633: Pixel = 145;
			7634: Pixel = 143;
			7635: Pixel = 142;
			7636: Pixel = 133;
			7637: Pixel = 123;
			7638: Pixel = 182;
			7639: Pixel = 218;
			7640: Pixel = 213;
			7641: Pixel = 212;
			7642: Pixel = 213;
			7643: Pixel = 216;
			7644: Pixel = 214;
			7645: Pixel = 210;
			7646: Pixel = 206;
			7647: Pixel = 205;
			7648: Pixel = 205;
			7649: Pixel = 205;
			7650: Pixel = 51;
			7651: Pixel = 52;
			7652: Pixel = 47;
			7653: Pixel = 59;
			7654: Pixel = 95;
			7655: Pixel = 107;
			7656: Pixel = 141;
			7657: Pixel = 162;
			7658: Pixel = 177;
			7659: Pixel = 178;
			7660: Pixel = 180;
			7661: Pixel = 166;
			7662: Pixel = 127;
			7663: Pixel = 68;
			7664: Pixel = 107;
			7665: Pixel = 111;
			7666: Pixel = 74;
			7667: Pixel = 73;
			7668: Pixel = 82;
			7669: Pixel = 41;
			7670: Pixel = 75;
			7671: Pixel = 46;
			7672: Pixel = 122;
			7673: Pixel = 128;
			7674: Pixel = 115;
			7675: Pixel = 118;
			7676: Pixel = 88;
			7677: Pixel = 121;
			7678: Pixel = 101;
			7679: Pixel = 104;
			7680: Pixel = 143;
			7681: Pixel = 199;
			7682: Pixel = 128;
			7683: Pixel = 40;
			7684: Pixel = 53;
			7685: Pixel = 53;
			7686: Pixel = 56;
			7687: Pixel = 50;
			7688: Pixel = 52;
			7689: Pixel = 54;
			7690: Pixel = 58;
			7691: Pixel = 60;
			7692: Pixel = 57;
			7693: Pixel = 59;
			7694: Pixel = 69;
			7695: Pixel = 66;
			7696: Pixel = 88;
			7697: Pixel = 102;
			7698: Pixel = 109;
			7699: Pixel = 121;
			7700: Pixel = 128;
			7701: Pixel = 133;
			7702: Pixel = 138;
			7703: Pixel = 138;
			7704: Pixel = 136;
			7705: Pixel = 134;
			7706: Pixel = 135;
			7707: Pixel = 138;
			7708: Pixel = 138;
			7709: Pixel = 140;
			7710: Pixel = 150;
			7711: Pixel = 150;
			7712: Pixel = 124;
			7713: Pixel = 59;
			7714: Pixel = 45;
			7715: Pixel = 45;
			7716: Pixel = 55;
			7717: Pixel = 59;
			7718: Pixel = 49;
			7719: Pixel = 63;
			7720: Pixel = 85;
			7721: Pixel = 76;
			7722: Pixel = 70;
			7723: Pixel = 63;
			7724: Pixel = 68;
			7725: Pixel = 160;
			7726: Pixel = 151;
			7727: Pixel = 150;
			7728: Pixel = 155;
			7729: Pixel = 154;
			7730: Pixel = 153;
			7731: Pixel = 153;
			7732: Pixel = 154;
			7733: Pixel = 152;
			7734: Pixel = 148;
			7735: Pixel = 146;
			7736: Pixel = 143;
			7737: Pixel = 141;
			7738: Pixel = 130;
			7739: Pixel = 119;
			7740: Pixel = 184;
			7741: Pixel = 221;
			7742: Pixel = 214;
			7743: Pixel = 214;
			7744: Pixel = 215;
			7745: Pixel = 215;
			7746: Pixel = 211;
			7747: Pixel = 207;
			7748: Pixel = 208;
			7749: Pixel = 209;
			7750: Pixel = 210;
			7751: Pixel = 210;
			7752: Pixel = 48;
			7753: Pixel = 50;
			7754: Pixel = 45;
			7755: Pixel = 68;
			7756: Pixel = 104;
			7757: Pixel = 112;
			7758: Pixel = 139;
			7759: Pixel = 161;
			7760: Pixel = 175;
			7761: Pixel = 176;
			7762: Pixel = 178;
			7763: Pixel = 166;
			7764: Pixel = 129;
			7765: Pixel = 72;
			7766: Pixel = 91;
			7767: Pixel = 110;
			7768: Pixel = 77;
			7769: Pixel = 86;
			7770: Pixel = 59;
			7771: Pixel = 46;
			7772: Pixel = 71;
			7773: Pixel = 49;
			7774: Pixel = 103;
			7775: Pixel = 114;
			7776: Pixel = 117;
			7777: Pixel = 130;
			7778: Pixel = 101;
			7779: Pixel = 89;
			7780: Pixel = 118;
			7781: Pixel = 97;
			7782: Pixel = 136;
			7783: Pixel = 172;
			7784: Pixel = 48;
			7785: Pixel = 50;
			7786: Pixel = 51;
			7787: Pixel = 54;
			7788: Pixel = 56;
			7789: Pixel = 49;
			7790: Pixel = 53;
			7791: Pixel = 49;
			7792: Pixel = 51;
			7793: Pixel = 58;
			7794: Pixel = 57;
			7795: Pixel = 53;
			7796: Pixel = 62;
			7797: Pixel = 60;
			7798: Pixel = 67;
			7799: Pixel = 85;
			7800: Pixel = 104;
			7801: Pixel = 115;
			7802: Pixel = 127;
			7803: Pixel = 133;
			7804: Pixel = 136;
			7805: Pixel = 139;
			7806: Pixel = 142;
			7807: Pixel = 150;
			7808: Pixel = 152;
			7809: Pixel = 164;
			7810: Pixel = 171;
			7811: Pixel = 163;
			7812: Pixel = 155;
			7813: Pixel = 153;
			7814: Pixel = 86;
			7815: Pixel = 48;
			7816: Pixel = 46;
			7817: Pixel = 50;
			7818: Pixel = 59;
			7819: Pixel = 58;
			7820: Pixel = 49;
			7821: Pixel = 67;
			7822: Pixel = 89;
			7823: Pixel = 78;
			7824: Pixel = 75;
			7825: Pixel = 66;
			7826: Pixel = 67;
			7827: Pixel = 162;
			7828: Pixel = 152;
			7829: Pixel = 152;
			7830: Pixel = 157;
			7831: Pixel = 154;
			7832: Pixel = 153;
			7833: Pixel = 151;
			7834: Pixel = 151;
			7835: Pixel = 151;
			7836: Pixel = 149;
			7837: Pixel = 145;
			7838: Pixel = 141;
			7839: Pixel = 139;
			7840: Pixel = 128;
			7841: Pixel = 119;
			7842: Pixel = 190;
			7843: Pixel = 222;
			7844: Pixel = 216;
			7845: Pixel = 213;
			7846: Pixel = 212;
			7847: Pixel = 212;
			7848: Pixel = 212;
			7849: Pixel = 212;
			7850: Pixel = 210;
			7851: Pixel = 208;
			7852: Pixel = 207;
			7853: Pixel = 206;
			7854: Pixel = 48;
			7855: Pixel = 49;
			7856: Pixel = 45;
			7857: Pixel = 70;
			7858: Pixel = 98;
			7859: Pixel = 112;
			7860: Pixel = 140;
			7861: Pixel = 162;
			7862: Pixel = 175;
			7863: Pixel = 176;
			7864: Pixel = 178;
			7865: Pixel = 166;
			7866: Pixel = 127;
			7867: Pixel = 74;
			7868: Pixel = 84;
			7869: Pixel = 95;
			7870: Pixel = 59;
			7871: Pixel = 85;
			7872: Pixel = 65;
			7873: Pixel = 51;
			7874: Pixel = 67;
			7875: Pixel = 48;
			7876: Pixel = 104;
			7877: Pixel = 87;
			7878: Pixel = 70;
			7879: Pixel = 124;
			7880: Pixel = 126;
			7881: Pixel = 106;
			7882: Pixel = 130;
			7883: Pixel = 113;
			7884: Pixel = 94;
			7885: Pixel = 90;
			7886: Pixel = 53;
			7887: Pixel = 53;
			7888: Pixel = 49;
			7889: Pixel = 58;
			7890: Pixel = 57;
			7891: Pixel = 50;
			7892: Pixel = 53;
			7893: Pixel = 52;
			7894: Pixel = 47;
			7895: Pixel = 53;
			7896: Pixel = 57;
			7897: Pixel = 55;
			7898: Pixel = 59;
			7899: Pixel = 61;
			7900: Pixel = 63;
			7901: Pixel = 50;
			7902: Pixel = 76;
			7903: Pixel = 99;
			7904: Pixel = 123;
			7905: Pixel = 132;
			7906: Pixel = 137;
			7907: Pixel = 144;
			7908: Pixel = 148;
			7909: Pixel = 159;
			7910: Pixel = 167;
			7911: Pixel = 167;
			7912: Pixel = 167;
			7913: Pixel = 171;
			7914: Pixel = 159;
			7915: Pixel = 143;
			7916: Pixel = 60;
			7917: Pixel = 54;
			7918: Pixel = 51;
			7919: Pixel = 53;
			7920: Pixel = 61;
			7921: Pixel = 54;
			7922: Pixel = 49;
			7923: Pixel = 73;
			7924: Pixel = 93;
			7925: Pixel = 79;
			7926: Pixel = 75;
			7927: Pixel = 67;
			7928: Pixel = 69;
			7929: Pixel = 162;
			7930: Pixel = 153;
			7931: Pixel = 153;
			7932: Pixel = 157;
			7933: Pixel = 152;
			7934: Pixel = 150;
			7935: Pixel = 150;
			7936: Pixel = 149;
			7937: Pixel = 150;
			7938: Pixel = 148;
			7939: Pixel = 143;
			7940: Pixel = 139;
			7941: Pixel = 137;
			7942: Pixel = 126;
			7943: Pixel = 124;
			7944: Pixel = 202;
			7945: Pixel = 222;
			7946: Pixel = 212;
			7947: Pixel = 210;
			7948: Pixel = 212;
			7949: Pixel = 214;
			7950: Pixel = 213;
			7951: Pixel = 207;
			7952: Pixel = 205;
			7953: Pixel = 207;
			7954: Pixel = 211;
			7955: Pixel = 201;
			7956: Pixel = 48;
			7957: Pixel = 48;
			7958: Pixel = 45;
			7959: Pixel = 57;
			7960: Pixel = 91;
			7961: Pixel = 117;
			7962: Pixel = 142;
			7963: Pixel = 163;
			7964: Pixel = 173;
			7965: Pixel = 175;
			7966: Pixel = 178;
			7967: Pixel = 167;
			7968: Pixel = 129;
			7969: Pixel = 59;
			7970: Pixel = 92;
			7971: Pixel = 84;
			7972: Pixel = 47;
			7973: Pixel = 84;
			7974: Pixel = 64;
			7975: Pixel = 61;
			7976: Pixel = 62;
			7977: Pixel = 39;
			7978: Pixel = 101;
			7979: Pixel = 115;
			7980: Pixel = 60;
			7981: Pixel = 96;
			7982: Pixel = 120;
			7983: Pixel = 129;
			7984: Pixel = 128;
			7985: Pixel = 137;
			7986: Pixel = 107;
			7987: Pixel = 72;
			7988: Pixel = 45;
			7989: Pixel = 54;
			7990: Pixel = 50;
			7991: Pixel = 60;
			7992: Pixel = 61;
			7993: Pixel = 52;
			7994: Pixel = 55;
			7995: Pixel = 53;
			7996: Pixel = 50;
			7997: Pixel = 49;
			7998: Pixel = 56;
			7999: Pixel = 57;
			8000: Pixel = 60;
			8001: Pixel = 59;
			8002: Pixel = 70;
			8003: Pixel = 56;
			8004: Pixel = 47;
			8005: Pixel = 67;
			8006: Pixel = 87;
			8007: Pixel = 101;
			8008: Pixel = 117;
			8009: Pixel = 129;
			8010: Pixel = 140;
			8011: Pixel = 148;
			8012: Pixel = 158;
			8013: Pixel = 168;
			8014: Pixel = 162;
			8015: Pixel = 159;
			8016: Pixel = 149;
			8017: Pixel = 120;
			8018: Pixel = 49;
			8019: Pixel = 57;
			8020: Pixel = 58;
			8021: Pixel = 55;
			8022: Pixel = 63;
			8023: Pixel = 55;
			8024: Pixel = 49;
			8025: Pixel = 78;
			8026: Pixel = 94;
			8027: Pixel = 79;
			8028: Pixel = 82;
			8029: Pixel = 73;
			8030: Pixel = 73;
			8031: Pixel = 160;
			8032: Pixel = 150;
			8033: Pixel = 138;
			8034: Pixel = 147;
			8035: Pixel = 148;
			8036: Pixel = 149;
			8037: Pixel = 151;
			8038: Pixel = 149;
			8039: Pixel = 149;
			8040: Pixel = 145;
			8041: Pixel = 141;
			8042: Pixel = 138;
			8043: Pixel = 136;
			8044: Pixel = 120;
			8045: Pixel = 134;
			8046: Pixel = 211;
			8047: Pixel = 220;
			8048: Pixel = 211;
			8049: Pixel = 211;
			8050: Pixel = 213;
			8051: Pixel = 213;
			8052: Pixel = 209;
			8053: Pixel = 206;
			8054: Pixel = 205;
			8055: Pixel = 183;
			8056: Pixel = 132;
			8057: Pixel = 87;
			8058: Pixel = 47;
			8059: Pixel = 47;
			8060: Pixel = 41;
			8061: Pixel = 49;
			8062: Pixel = 84;
			8063: Pixel = 103;
			8064: Pixel = 141;
			8065: Pixel = 164;
			8066: Pixel = 173;
			8067: Pixel = 173;
			8068: Pixel = 176;
			8069: Pixel = 166;
			8070: Pixel = 110;
			8071: Pixel = 107;
			8072: Pixel = 137;
			8073: Pixel = 101;
			8074: Pixel = 54;
			8075: Pixel = 72;
			8076: Pixel = 61;
			8077: Pixel = 63;
			8078: Pixel = 53;
			8079: Pixel = 38;
			8080: Pixel = 85;
			8081: Pixel = 143;
			8082: Pixel = 87;
			8083: Pixel = 72;
			8084: Pixel = 105;
			8085: Pixel = 100;
			8086: Pixel = 126;
			8087: Pixel = 147;
			8088: Pixel = 124;
			8089: Pixel = 136;
			8090: Pixel = 59;
			8091: Pixel = 42;
			8092: Pixel = 50;
			8093: Pixel = 69;
			8094: Pixel = 61;
			8095: Pixel = 50;
			8096: Pixel = 55;
			8097: Pixel = 49;
			8098: Pixel = 51;
			8099: Pixel = 48;
			8100: Pixel = 51;
			8101: Pixel = 59;
			8102: Pixel = 61;
			8103: Pixel = 58;
			8104: Pixel = 62;
			8105: Pixel = 76;
			8106: Pixel = 72;
			8107: Pixel = 87;
			8108: Pixel = 97;
			8109: Pixel = 111;
			8110: Pixel = 119;
			8111: Pixel = 126;
			8112: Pixel = 135;
			8113: Pixel = 149;
			8114: Pixel = 154;
			8115: Pixel = 161;
			8116: Pixel = 162;
			8117: Pixel = 157;
			8118: Pixel = 153;
			8119: Pixel = 136;
			8120: Pixel = 66;
			8121: Pixel = 47;
			8122: Pixel = 51;
			8123: Pixel = 57;
			8124: Pixel = 62;
			8125: Pixel = 53;
			8126: Pixel = 50;
			8127: Pixel = 77;
			8128: Pixel = 96;
			8129: Pixel = 83;
			8130: Pixel = 84;
			8131: Pixel = 71;
			8132: Pixel = 82;
			8133: Pixel = 162;
			8134: Pixel = 132;
			8135: Pixel = 111;
			8136: Pixel = 121;
			8137: Pixel = 130;
			8138: Pixel = 134;
			8139: Pixel = 139;
			8140: Pixel = 144;
			8141: Pixel = 148;
			8142: Pixel = 146;
			8143: Pixel = 142;
			8144: Pixel = 137;
			8145: Pixel = 132;
			8146: Pixel = 114;
			8147: Pixel = 152;
			8148: Pixel = 218;
			8149: Pixel = 214;
			8150: Pixel = 210;
			8151: Pixel = 210;
			8152: Pixel = 209;
			8153: Pixel = 208;
			8154: Pixel = 201;
			8155: Pixel = 185;
			8156: Pixel = 128;
			8157: Pixel = 63;
			8158: Pixel = 34;
			8159: Pixel = 42;
			8160: Pixel = 56;
			8161: Pixel = 54;
			8162: Pixel = 42;
			8163: Pixel = 47;
			8164: Pixel = 70;
			8165: Pixel = 90;
			8166: Pixel = 138;
			8167: Pixel = 162;
			8168: Pixel = 173;
			8169: Pixel = 172;
			8170: Pixel = 175;
			8171: Pixel = 156;
			8172: Pixel = 147;
			8173: Pixel = 146;
			8174: Pixel = 75;
			8175: Pixel = 87;
			8176: Pixel = 41;
			8177: Pixel = 76;
			8178: Pixel = 66;
			8179: Pixel = 60;
			8180: Pixel = 68;
			8181: Pixel = 47;
			8182: Pixel = 78;
			8183: Pixel = 132;
			8184: Pixel = 117;
			8185: Pixel = 59;
			8186: Pixel = 91;
			8187: Pixel = 134;
			8188: Pixel = 95;
			8189: Pixel = 130;
			8190: Pixel = 91;
			8191: Pixel = 106;
			8192: Pixel = 153;
			8193: Pixel = 57;
			8194: Pixel = 44;
			8195: Pixel = 73;
			8196: Pixel = 60;
			8197: Pixel = 55;
			8198: Pixel = 56;
			8199: Pixel = 49;
			8200: Pixel = 52;
			8201: Pixel = 49;
			8202: Pixel = 51;
			8203: Pixel = 56;
			8204: Pixel = 59;
			8205: Pixel = 54;
			8206: Pixel = 52;
			8207: Pixel = 79;
			8208: Pixel = 105;
			8209: Pixel = 129;
			8210: Pixel = 132;
			8211: Pixel = 134;
			8212: Pixel = 137;
			8213: Pixel = 137;
			8214: Pixel = 142;
			8215: Pixel = 150;
			8216: Pixel = 151;
			8217: Pixel = 149;
			8218: Pixel = 151;
			8219: Pixel = 162;
			8220: Pixel = 181;
			8221: Pixel = 198;
			8222: Pixel = 189;
			8223: Pixel = 142;
			8224: Pixel = 80;
			8225: Pixel = 46;
			8226: Pixel = 49;
			8227: Pixel = 52;
			8228: Pixel = 51;
			8229: Pixel = 80;
			8230: Pixel = 93;
			8231: Pixel = 82;
			8232: Pixel = 83;
			8233: Pixel = 74;
			8234: Pixel = 89;
			8235: Pixel = 159;
			8236: Pixel = 121;
			8237: Pixel = 116;
			8238: Pixel = 112;
			8239: Pixel = 113;
			8240: Pixel = 113;
			8241: Pixel = 114;
			8242: Pixel = 119;
			8243: Pixel = 128;
			8244: Pixel = 133;
			8245: Pixel = 134;
			8246: Pixel = 135;
			8247: Pixel = 129;
			8248: Pixel = 114;
			8249: Pixel = 170;
			8250: Pixel = 219;
			8251: Pixel = 207;
			8252: Pixel = 207;
			8253: Pixel = 209;
			8254: Pixel = 206;
			8255: Pixel = 200;
			8256: Pixel = 191;
			8257: Pixel = 128;
			8258: Pixel = 44;
			8259: Pixel = 38;
			8260: Pixel = 63;
			8261: Pixel = 78;
			8262: Pixel = 98;
			8263: Pixel = 74;
			8264: Pixel = 55;
			8265: Pixel = 53;
			8266: Pixel = 60;
			8267: Pixel = 69;
			8268: Pixel = 123;
			8269: Pixel = 160;
			8270: Pixel = 171;
			8271: Pixel = 170;
			8272: Pixel = 174;
			8273: Pixel = 175;
			8274: Pixel = 152;
			8275: Pixel = 64;
			8276: Pixel = 101;
			8277: Pixel = 78;
			8278: Pixel = 31;
			8279: Pixel = 63;
			8280: Pixel = 68;
			8281: Pixel = 48;
			8282: Pixel = 79;
			8283: Pixel = 77;
			8284: Pixel = 54;
			8285: Pixel = 95;
			8286: Pixel = 120;
			8287: Pixel = 92;
			8288: Pixel = 130;
			8289: Pixel = 112;
			8290: Pixel = 83;
			8291: Pixel = 108;
			8292: Pixel = 102;
			8293: Pixel = 122;
			8294: Pixel = 128;
			8295: Pixel = 111;
			8296: Pixel = 48;
			8297: Pixel = 69;
			8298: Pixel = 55;
			8299: Pixel = 58;
			8300: Pixel = 59;
			8301: Pixel = 47;
			8302: Pixel = 51;
			8303: Pixel = 52;
			8304: Pixel = 49;
			8305: Pixel = 53;
			8306: Pixel = 61;
			8307: Pixel = 57;
			8308: Pixel = 52;
			8309: Pixel = 77;
			8310: Pixel = 111;
			8311: Pixel = 124;
			8312: Pixel = 124;
			8313: Pixel = 124;
			8314: Pixel = 132;
			8315: Pixel = 136;
			8316: Pixel = 138;
			8317: Pixel = 143;
			8318: Pixel = 141;
			8319: Pixel = 141;
			8320: Pixel = 145;
			8321: Pixel = 163;
			8322: Pixel = 182;
			8323: Pixel = 194;
			8324: Pixel = 202;
			8325: Pixel = 211;
			8326: Pixel = 200;
			8327: Pixel = 150;
			8328: Pixel = 73;
			8329: Pixel = 33;
			8330: Pixel = 43;
			8331: Pixel = 82;
			8332: Pixel = 89;
			8333: Pixel = 78;
			8334: Pixel = 80;
			8335: Pixel = 69;
			8336: Pixel = 95;
			8337: Pixel = 155;
			8338: Pixel = 128;
			8339: Pixel = 135;
			8340: Pixel = 130;
			8341: Pixel = 122;
			8342: Pixel = 115;
			8343: Pixel = 107;
			8344: Pixel = 102;
			8345: Pixel = 101;
			8346: Pixel = 105;
			8347: Pixel = 107;
			8348: Pixel = 110;
			8349: Pixel = 113;
			8350: Pixel = 101;
			8351: Pixel = 167;
			8352: Pixel = 213;
			8353: Pixel = 203;
			8354: Pixel = 207;
			8355: Pixel = 208;
			8356: Pixel = 208;
			8357: Pixel = 194;
			8358: Pixel = 127;
			8359: Pixel = 53;
			8360: Pixel = 50;
			8361: Pixel = 67;
			8362: Pixel = 83;
			8363: Pixel = 86;
			8364: Pixel = 136;
			8365: Pixel = 121;
			8366: Pixel = 88;
			8367: Pixel = 73;
			8368: Pixel = 58;
			8369: Pixel = 55;
			8370: Pixel = 113;
			8371: Pixel = 159;
			8372: Pixel = 169;
			8373: Pixel = 169;
			8374: Pixel = 175;
			8375: Pixel = 173;
			8376: Pixel = 116;
			8377: Pixel = 107;
			8378: Pixel = 129;
			8379: Pixel = 38;
			8380: Pixel = 40;
			8381: Pixel = 47;
			8382: Pixel = 97;
			8383: Pixel = 37;
			8384: Pixel = 76;
			8385: Pixel = 101;
			8386: Pixel = 65;
			8387: Pixel = 45;
			8388: Pixel = 110;
			8389: Pixel = 102;
			8390: Pixel = 109;
			8391: Pixel = 80;
			8392: Pixel = 107;
			8393: Pixel = 109;
			8394: Pixel = 122;
			8395: Pixel = 131;
			8396: Pixel = 109;
			8397: Pixel = 84;
			8398: Pixel = 92;
			8399: Pixel = 58;
			8400: Pixel = 52;
			8401: Pixel = 58;
			8402: Pixel = 59;
			8403: Pixel = 48;
			8404: Pixel = 49;
			8405: Pixel = 58;
			8406: Pixel = 50;
			8407: Pixel = 52;
			8408: Pixel = 60;
			8409: Pixel = 66;
			8410: Pixel = 50;
			8411: Pixel = 72;
			8412: Pixel = 108;
			8413: Pixel = 118;
			8414: Pixel = 123;
			8415: Pixel = 127;
			8416: Pixel = 129;
			8417: Pixel = 137;
			8418: Pixel = 139;
			8419: Pixel = 139;
			8420: Pixel = 139;
			8421: Pixel = 143;
			8422: Pixel = 153;
			8423: Pixel = 169;
			8424: Pixel = 185;
			8425: Pixel = 190;
			8426: Pixel = 193;
			8427: Pixel = 196;
			8428: Pixel = 202;
			8429: Pixel = 215;
			8430: Pixel = 204;
			8431: Pixel = 110;
			8432: Pixel = 33;
			8433: Pixel = 70;
			8434: Pixel = 86;
			8435: Pixel = 74;
			8436: Pixel = 76;
			8437: Pixel = 64;
			8438: Pixel = 99;
			8439: Pixel = 153;
			8440: Pixel = 140;
			8441: Pixel = 142;
			8442: Pixel = 140;
			8443: Pixel = 134;
			8444: Pixel = 132;
			8445: Pixel = 125;
			8446: Pixel = 115;
			8447: Pixel = 106;
			8448: Pixel = 98;
			8449: Pixel = 90;
			8450: Pixel = 101;
			8451: Pixel = 116;
			8452: Pixel = 77;
			8453: Pixel = 153;
			8454: Pixel = 212;
			8455: Pixel = 205;
			8456: Pixel = 209;
			8457: Pixel = 206;
			8458: Pixel = 195;
			8459: Pixel = 130;
			8460: Pixel = 48;
			8461: Pixel = 65;
			8462: Pixel = 76;
			8463: Pixel = 80;
			8464: Pixel = 86;
			8465: Pixel = 85;
			8466: Pixel = 134;
			8467: Pixel = 145;
			8468: Pixel = 131;
			8469: Pixel = 102;
			8470: Pixel = 66;
			8471: Pixel = 51;
			8472: Pixel = 114;
			8473: Pixel = 160;
			8474: Pixel = 171;
			8475: Pixel = 170;
			8476: Pixel = 174;
			8477: Pixel = 158;
			8478: Pixel = 149;
			8479: Pixel = 145;
			8480: Pixel = 76;
			8481: Pixel = 42;
			8482: Pixel = 38;
			8483: Pixel = 49;
			8484: Pixel = 96;
			8485: Pixel = 92;
			8486: Pixel = 99;
			8487: Pixel = 75;
			8488: Pixel = 71;
			8489: Pixel = 84;
			8490: Pixel = 68;
			8491: Pixel = 104;
			8492: Pixel = 75;
			8493: Pixel = 70;
			8494: Pixel = 98;
			8495: Pixel = 121;
			8496: Pixel = 142;
			8497: Pixel = 124;
			8498: Pixel = 88;
			8499: Pixel = 87;
			8500: Pixel = 104;
			8501: Pixel = 69;
			8502: Pixel = 44;
			8503: Pixel = 62;
			8504: Pixel = 62;
			8505: Pixel = 52;
			8506: Pixel = 49;
			8507: Pixel = 60;
			8508: Pixel = 56;
			8509: Pixel = 52;
			8510: Pixel = 61;
			8511: Pixel = 75;
			8512: Pixel = 55;
			8513: Pixel = 71;
			8514: Pixel = 107;
			8515: Pixel = 119;
			8516: Pixel = 124;
			8517: Pixel = 124;
			8518: Pixel = 133;
			8519: Pixel = 140;
			8520: Pixel = 142;
			8521: Pixel = 137;
			8522: Pixel = 138;
			8523: Pixel = 148;
			8524: Pixel = 158;
			8525: Pixel = 168;
			8526: Pixel = 180;
			8527: Pixel = 186;
			8528: Pixel = 189;
			8529: Pixel = 193;
			8530: Pixel = 199;
			8531: Pixel = 201;
			8532: Pixel = 210;
			8533: Pixel = 222;
			8534: Pixel = 135;
			8535: Pixel = 46;
			8536: Pixel = 76;
			8537: Pixel = 65;
			8538: Pixel = 76;
			8539: Pixel = 57;
			8540: Pixel = 104;
			8541: Pixel = 152;
			8542: Pixel = 145;
			8543: Pixel = 147;
			8544: Pixel = 143;
			8545: Pixel = 141;
			8546: Pixel = 139;
			8547: Pixel = 135;
			8548: Pixel = 130;
			8549: Pixel = 122;
			8550: Pixel = 116;
			8551: Pixel = 103;
			8552: Pixel = 116;
			8553: Pixel = 128;
			8554: Pixel = 88;
			8555: Pixel = 172;
			8556: Pixel = 215;
			8557: Pixel = 210;
			8558: Pixel = 210;
			8559: Pixel = 208;
			8560: Pixel = 133;
			8561: Pixel = 41;
			8562: Pixel = 74;
			8563: Pixel = 86;
			8564: Pixel = 80;
			8565: Pixel = 95;
			8566: Pixel = 92;
			8567: Pixel = 84;
			8568: Pixel = 127;
			8569: Pixel = 146;
			8570: Pixel = 150;
			8571: Pixel = 133;
			8572: Pixel = 82;
			8573: Pixel = 50;
			8574: Pixel = 113;
			8575: Pixel = 162;
			8576: Pixel = 175;
			8577: Pixel = 173;
			8578: Pixel = 177;
			8579: Pixel = 156;
			8580: Pixel = 173;
			8581: Pixel = 145;
			8582: Pixel = 63;
			8583: Pixel = 45;
			8584: Pixel = 51;
			8585: Pixel = 59;
			8586: Pixel = 55;
			8587: Pixel = 68;
			8588: Pixel = 62;
			8589: Pixel = 59;
			8590: Pixel = 67;
			8591: Pixel = 62;
			8592: Pixel = 65;
			8593: Pixel = 93;
			8594: Pixel = 54;
			8595: Pixel = 75;
			8596: Pixel = 93;
			8597: Pixel = 103;
			8598: Pixel = 137;
			8599: Pixel = 141;
			8600: Pixel = 83;
			8601: Pixel = 127;
			8602: Pixel = 107;
			8603: Pixel = 85;
			8604: Pixel = 39;
			8605: Pixel = 63;
			8606: Pixel = 62;
			8607: Pixel = 54;
			8608: Pixel = 52;
			8609: Pixel = 62;
			8610: Pixel = 57;
			8611: Pixel = 57;
			8612: Pixel = 66;
			8613: Pixel = 92;
			8614: Pixel = 68;
			8615: Pixel = 60;
			8616: Pixel = 114;
			8617: Pixel = 121;
			8618: Pixel = 118;
			8619: Pixel = 130;
			8620: Pixel = 138;
			8621: Pixel = 137;
			8622: Pixel = 140;
			8623: Pixel = 139;
			8624: Pixel = 143;
			8625: Pixel = 153;
			8626: Pixel = 161;
			8627: Pixel = 166;
			8628: Pixel = 173;
			8629: Pixel = 179;
			8630: Pixel = 184;
			8631: Pixel = 189;
			8632: Pixel = 194;
			8633: Pixel = 201;
			8634: Pixel = 205;
			8635: Pixel = 209;
			8636: Pixel = 226;
			8637: Pixel = 131;
			8638: Pixel = 49;
			8639: Pixel = 58;
			8640: Pixel = 75;
			8641: Pixel = 55;
			8642: Pixel = 111;
			8643: Pixel = 151;
			8644: Pixel = 145;
			8645: Pixel = 147;
			8646: Pixel = 143;
			8647: Pixel = 143;
			8648: Pixel = 141;
			8649: Pixel = 138;
			8650: Pixel = 135;
			8651: Pixel = 130;
			8652: Pixel = 127;
			8653: Pixel = 119;
			8654: Pixel = 123;
			8655: Pixel = 126;
			8656: Pixel = 120;
			8657: Pixel = 197;
			8658: Pixel = 213;
			8659: Pixel = 212;
			8660: Pixel = 209;
			8661: Pixel = 186;
			8662: Pixel = 84;
			8663: Pixel = 61;
			8664: Pixel = 96;
			8665: Pixel = 87;
			8666: Pixel = 96;
			8667: Pixel = 108;
			8668: Pixel = 91;
			8669: Pixel = 92;
			8670: Pixel = 84;
			8671: Pixel = 131;
			8672: Pixel = 157;
			8673: Pixel = 158;
			8674: Pixel = 103;
			8675: Pixel = 49;
			8676: Pixel = 113;
			8677: Pixel = 163;
			8678: Pixel = 176;
			8679: Pixel = 176;
			8680: Pixel = 179;
			8681: Pixel = 160;
			8682: Pixel = 160;
			8683: Pixel = 111;
			8684: Pixel = 48;
			8685: Pixel = 40;
			8686: Pixel = 47;
			8687: Pixel = 62;
			8688: Pixel = 60;
			8689: Pixel = 43;
			8690: Pixel = 62;
			8691: Pixel = 83;
			8692: Pixel = 42;
			8693: Pixel = 58;
			8694: Pixel = 57;
			8695: Pixel = 78;
			8696: Pixel = 71;
			8697: Pixel = 67;
			8698: Pixel = 82;
			8699: Pixel = 101;
			8700: Pixel = 126;
			8701: Pixel = 128;
			8702: Pixel = 136;
			8703: Pixel = 99;
			8704: Pixel = 113;
			8705: Pixel = 110;
			8706: Pixel = 36;
			8707: Pixel = 59;
			8708: Pixel = 63;
			8709: Pixel = 52;
			8710: Pixel = 47;
			8711: Pixel = 61;
			8712: Pixel = 57;
			8713: Pixel = 50;
			8714: Pixel = 64;
			8715: Pixel = 107;
			8716: Pixel = 85;
			8717: Pixel = 54;
			8718: Pixel = 110;
			8719: Pixel = 118;
			8720: Pixel = 130;
			8721: Pixel = 134;
			8722: Pixel = 138;
			8723: Pixel = 139;
			8724: Pixel = 138;
			8725: Pixel = 140;
			8726: Pixel = 145;
			8727: Pixel = 152;
			8728: Pixel = 159;
			8729: Pixel = 162;
			8730: Pixel = 169;
			8731: Pixel = 174;
			8732: Pixel = 179;
			8733: Pixel = 184;
			8734: Pixel = 192;
			8735: Pixel = 198;
			8736: Pixel = 204;
			8737: Pixel = 208;
			8738: Pixel = 214;
			8739: Pixel = 223;
			8740: Pixel = 94;
			8741: Pixel = 39;
			8742: Pixel = 65;
			8743: Pixel = 49;
			8744: Pixel = 121;
			8745: Pixel = 147;
			8746: Pixel = 146;
			8747: Pixel = 146;
			8748: Pixel = 143;
			8749: Pixel = 143;
			8750: Pixel = 142;
			8751: Pixel = 141;
			8752: Pixel = 136;
			8753: Pixel = 134;
			8754: Pixel = 129;
			8755: Pixel = 125;
			8756: Pixel = 131;
			8757: Pixel = 129;
			8758: Pixel = 144;
			8759: Pixel = 210;
			8760: Pixel = 213;
			8761: Pixel = 212;
			8762: Pixel = 207;
			8763: Pixel = 145;
			8764: Pixel = 72;
			8765: Pixel = 91;
			8766: Pixel = 92;
			8767: Pixel = 96;
			8768: Pixel = 112;
			8769: Pixel = 103;
			8770: Pixel = 92;
			8771: Pixel = 101;
			8772: Pixel = 42;
			8773: Pixel = 105;
			8774: Pixel = 164;
			8775: Pixel = 167;
			8776: Pixel = 121;
			8777: Pixel = 46;
			8778: Pixel = 109;
			8779: Pixel = 165;
			8780: Pixel = 176;
			8781: Pixel = 176;
			8782: Pixel = 178;
			8783: Pixel = 162;
			8784: Pixel = 150;
			8785: Pixel = 115;
			8786: Pixel = 44;
			8787: Pixel = 41;
			8788: Pixel = 52;
			8789: Pixel = 62;
			8790: Pixel = 48;
			8791: Pixel = 44;
			8792: Pixel = 76;
			8793: Pixel = 83;
			8794: Pixel = 54;
			8795: Pixel = 47;
			8796: Pixel = 71;
			8797: Pixel = 68;
			8798: Pixel = 78;
			8799: Pixel = 86;
			8800: Pixel = 89;
			8801: Pixel = 87;
			8802: Pixel = 106;
			8803: Pixel = 125;
			8804: Pixel = 158;
			8805: Pixel = 69;
			8806: Pixel = 85;
			8807: Pixel = 151;
			8808: Pixel = 39;
			8809: Pixel = 51;
			8810: Pixel = 65;
			8811: Pixel = 51;
			8812: Pixel = 45;
			8813: Pixel = 61;
			8814: Pixel = 58;
			8815: Pixel = 48;
			8816: Pixel = 62;
			8817: Pixel = 116;
			8818: Pixel = 91;
			8819: Pixel = 49;
			8820: Pixel = 104;
			8821: Pixel = 127;
			8822: Pixel = 133;
			8823: Pixel = 132;
			8824: Pixel = 136;
			8825: Pixel = 140;
			8826: Pixel = 140;
			8827: Pixel = 141;
			8828: Pixel = 146;
			8829: Pixel = 150;
			8830: Pixel = 155;
			8831: Pixel = 161;
			8832: Pixel = 165;
			8833: Pixel = 171;
			8834: Pixel = 177;
			8835: Pixel = 183;
			8836: Pixel = 190;
			8837: Pixel = 196;
			8838: Pixel = 202;
			8839: Pixel = 207;
			8840: Pixel = 209;
			8841: Pixel = 226;
			8842: Pixel = 191;
			8843: Pixel = 47;
			8844: Pixel = 51;
			8845: Pixel = 46;
			8846: Pixel = 128;
			8847: Pixel = 144;
			8848: Pixel = 146;
			8849: Pixel = 145;
			8850: Pixel = 144;
			8851: Pixel = 142;
			8852: Pixel = 140;
			8853: Pixel = 139;
			8854: Pixel = 138;
			8855: Pixel = 136;
			8856: Pixel = 130;
			8857: Pixel = 125;
			8858: Pixel = 128;
			8859: Pixel = 145;
			8860: Pixel = 173;
			8861: Pixel = 214;
			8862: Pixel = 213;
			8863: Pixel = 212;
			8864: Pixel = 197;
			8865: Pixel = 104;
			8866: Pixel = 80;
			8867: Pixel = 93;
			8868: Pixel = 98;
			8869: Pixel = 110;
			8870: Pixel = 103;
			8871: Pixel = 89;
			8872: Pixel = 101;
			8873: Pixel = 104;
			8874: Pixel = 33;
			8875: Pixel = 84;
			8876: Pixel = 164;
			8877: Pixel = 173;
			8878: Pixel = 125;
			8879: Pixel = 38;
			8880: Pixel = 107;
			8881: Pixel = 164;
			8882: Pixel = 177;
			8883: Pixel = 176;
			8884: Pixel = 179;
			8885: Pixel = 169;
			8886: Pixel = 135;
			8887: Pixel = 112;
			8888: Pixel = 48;
			8889: Pixel = 44;
			8890: Pixel = 57;
			8891: Pixel = 49;
			8892: Pixel = 49;
			8893: Pixel = 40;
			8894: Pixel = 89;
			8895: Pixel = 77;
			8896: Pixel = 58;
			8897: Pixel = 42;
			8898: Pixel = 56;
			8899: Pixel = 78;
			8900: Pixel = 64;
			8901: Pixel = 84;
			8902: Pixel = 108;
			8903: Pixel = 85;
			8904: Pixel = 92;
			8905: Pixel = 143;
			8906: Pixel = 144;
			8907: Pixel = 55;
			8908: Pixel = 86;
			8909: Pixel = 165;
			8910: Pixel = 33;
			8911: Pixel = 55;
			8912: Pixel = 72;
			8913: Pixel = 55;
			8914: Pixel = 47;
			8915: Pixel = 60;
			8916: Pixel = 52;
			8917: Pixel = 48;
			8918: Pixel = 74;
			8919: Pixel = 110;
			8920: Pixel = 90;
			8921: Pixel = 54;
			8922: Pixel = 107;
			8923: Pixel = 128;
			8924: Pixel = 128;
			8925: Pixel = 134;
			8926: Pixel = 137;
			8927: Pixel = 138;
			8928: Pixel = 140;
			8929: Pixel = 142;
			8930: Pixel = 147;
			8931: Pixel = 148;
			8932: Pixel = 153;
			8933: Pixel = 158;
			8934: Pixel = 163;
			8935: Pixel = 170;
			8936: Pixel = 175;
			8937: Pixel = 182;
			8938: Pixel = 187;
			8939: Pixel = 194;
			8940: Pixel = 202;
			8941: Pixel = 208;
			8942: Pixel = 211;
			8943: Pixel = 214;
			8944: Pixel = 231;
			8945: Pixel = 106;
			8946: Pixel = 28;
			8947: Pixel = 47;
			8948: Pixel = 138;
			8949: Pixel = 146;
			8950: Pixel = 149;
			8951: Pixel = 145;
			8952: Pixel = 144;
			8953: Pixel = 142;
			8954: Pixel = 140;
			8955: Pixel = 136;
			8956: Pixel = 135;
			8957: Pixel = 133;
			8958: Pixel = 127;
			8959: Pixel = 120;
			8960: Pixel = 149;
			8961: Pixel = 187;
			8962: Pixel = 203;
			8963: Pixel = 214;
			8964: Pixel = 213;
			8965: Pixel = 212;
			8966: Pixel = 166;
			8967: Pixel = 89;
			8968: Pixel = 93;
			8969: Pixel = 95;
			8970: Pixel = 108;
			8971: Pixel = 110;
			8972: Pixel = 90;
			8973: Pixel = 93;
			8974: Pixel = 103;
			8975: Pixel = 101;
			8976: Pixel = 31;
			8977: Pixel = 75;
			8978: Pixel = 157;
			8979: Pixel = 175;
			8980: Pixel = 122;
			8981: Pixel = 36;
			8982: Pixel = 105;
			8983: Pixel = 165;
			8984: Pixel = 178;
			8985: Pixel = 177;
			8986: Pixel = 181;
			8987: Pixel = 167;
			8988: Pixel = 150;
			8989: Pixel = 108;
			8990: Pixel = 43;
			8991: Pixel = 53;
			8992: Pixel = 52;
			8993: Pixel = 46;
			8994: Pixel = 47;
			8995: Pixel = 40;
			8996: Pixel = 119;
			8997: Pixel = 68;
			8998: Pixel = 47;
			8999: Pixel = 57;
			9000: Pixel = 55;
			9001: Pixel = 48;
			9002: Pixel = 53;
			9003: Pixel = 75;
			9004: Pixel = 103;
			9005: Pixel = 84;
			9006: Pixel = 81;
			9007: Pixel = 136;
			9008: Pixel = 142;
			9009: Pixel = 84;
			9010: Pixel = 84;
			9011: Pixel = 147;
			9012: Pixel = 43;
			9013: Pixel = 62;
			9014: Pixel = 72;
			9015: Pixel = 56;
			9016: Pixel = 49;
			9017: Pixel = 56;
			9018: Pixel = 52;
			9019: Pixel = 51;
			9020: Pixel = 85;
			9021: Pixel = 116;
			9022: Pixel = 102;
			9023: Pixel = 58;
			9024: Pixel = 108;
			9025: Pixel = 131;
			9026: Pixel = 131;
			9027: Pixel = 136;
			9028: Pixel = 138;
			9029: Pixel = 136;
			9030: Pixel = 137;
			9031: Pixel = 140;
			9032: Pixel = 145;
			9033: Pixel = 146;
			9034: Pixel = 152;
			9035: Pixel = 155;
			9036: Pixel = 162;
			9037: Pixel = 167;
			9038: Pixel = 173;
			9039: Pixel = 180;
			9040: Pixel = 186;
			9041: Pixel = 193;
			9042: Pixel = 201;
			9043: Pixel = 207;
			9044: Pixel = 210;
			9045: Pixel = 212;
			9046: Pixel = 228;
			9047: Pixel = 177;
			9048: Pixel = 27;
			9049: Pixel = 51;
			9050: Pixel = 143;
			9051: Pixel = 147;
			9052: Pixel = 148;
			9053: Pixel = 146;
			9054: Pixel = 145;
			9055: Pixel = 142;
			9056: Pixel = 139;
			9057: Pixel = 134;
			9058: Pixel = 133;
			9059: Pixel = 129;
			9060: Pixel = 122;
			9061: Pixel = 134;
			9062: Pixel = 198;
			9063: Pixel = 207;
			9064: Pixel = 206;
			9065: Pixel = 216;
			9066: Pixel = 215;
			9067: Pixel = 201;
			9068: Pixel = 126;
			9069: Pixel = 87;
			9070: Pixel = 93;
			9071: Pixel = 104;
			9072: Pixel = 115;
			9073: Pixel = 100;
			9074: Pixel = 89;
			9075: Pixel = 102;
			9076: Pixel = 101;
			9077: Pixel = 102;
			9078: Pixel = 27;
			9079: Pixel = 62;
			9080: Pixel = 153;
			9081: Pixel = 176;
			9082: Pixel = 130;
			9083: Pixel = 37;
			9084: Pixel = 101;
			9085: Pixel = 166;
			9086: Pixel = 178;
			9087: Pixel = 178;
			9088: Pixel = 181;
			9089: Pixel = 168;
			9090: Pixel = 147;
			9091: Pixel = 79;
			9092: Pixel = 49;
			9093: Pixel = 52;
			9094: Pixel = 43;
			9095: Pixel = 45;
			9096: Pixel = 38;
			9097: Pixel = 75;
			9098: Pixel = 112;
			9099: Pixel = 56;
			9100: Pixel = 42;
			9101: Pixel = 63;
			9102: Pixel = 48;
			9103: Pixel = 46;
			9104: Pixel = 53;
			9105: Pixel = 55;
			9106: Pixel = 94;
			9107: Pixel = 96;
			9108: Pixel = 80;
			9109: Pixel = 144;
			9110: Pixel = 136;
			9111: Pixel = 120;
			9112: Pixel = 140;
			9113: Pixel = 119;
			9114: Pixel = 61;
			9115: Pixel = 54;
			9116: Pixel = 60;
			9117: Pixel = 57;
			9118: Pixel = 55;
			9119: Pixel = 51;
			9120: Pixel = 52;
			9121: Pixel = 66;
			9122: Pixel = 109;
			9123: Pixel = 130;
			9124: Pixel = 100;
			9125: Pixel = 65;
			9126: Pixel = 112;
			9127: Pixel = 130;
			9128: Pixel = 135;
			9129: Pixel = 137;
			9130: Pixel = 136;
			9131: Pixel = 136;
			9132: Pixel = 137;
			9133: Pixel = 139;
			9134: Pixel = 143;
			9135: Pixel = 146;
			9136: Pixel = 149;
			9137: Pixel = 155;
			9138: Pixel = 160;
			9139: Pixel = 163;
			9140: Pixel = 172;
			9141: Pixel = 178;
			9142: Pixel = 185;
			9143: Pixel = 192;
			9144: Pixel = 199;
			9145: Pixel = 207;
			9146: Pixel = 210;
			9147: Pixel = 212;
			9148: Pixel = 217;
			9149: Pixel = 219;
			9150: Pixel = 54;
			9151: Pixel = 53;
			9152: Pixel = 146;
			9153: Pixel = 148;
			9154: Pixel = 146;
			9155: Pixel = 144;
			9156: Pixel = 143;
			9157: Pixel = 140;
			9158: Pixel = 139;
			9159: Pixel = 135;
			9160: Pixel = 131;
			9161: Pixel = 127;
			9162: Pixel = 118;
			9163: Pixel = 154;
			9164: Pixel = 219;
			9165: Pixel = 212;
			9166: Pixel = 210;
			9167: Pixel = 216;
			9168: Pixel = 215;
			9169: Pixel = 173;
			9170: Pixel = 104;
			9171: Pixel = 92;
			9172: Pixel = 93;
			9173: Pixel = 110;
			9174: Pixel = 111;
			9175: Pixel = 93;
			9176: Pixel = 96;
			9177: Pixel = 105;
			9178: Pixel = 101;
			9179: Pixel = 94;
			9180: Pixel = 27;
			9181: Pixel = 59;
			9182: Pixel = 150;
			9183: Pixel = 175;
			9184: Pixel = 137;
			9185: Pixel = 45;
			9186: Pixel = 97;
			9187: Pixel = 166;
			9188: Pixel = 176;
			9189: Pixel = 173;
			9190: Pixel = 175;
			9191: Pixel = 166;
			9192: Pixel = 143;
			9193: Pixel = 90;
			9194: Pixel = 51;
			9195: Pixel = 44;
			9196: Pixel = 46;
			9197: Pixel = 48;
			9198: Pixel = 65;
			9199: Pixel = 62;
			9200: Pixel = 81;
			9201: Pixel = 65;
			9202: Pixel = 47;
			9203: Pixel = 64;
			9204: Pixel = 43;
			9205: Pixel = 49;
			9206: Pixel = 55;
			9207: Pixel = 66;
			9208: Pixel = 59;
			9209: Pixel = 91;
			9210: Pixel = 129;
			9211: Pixel = 136;
			9212: Pixel = 102;
			9213: Pixel = 117;
			9214: Pixel = 152;
			9215: Pixel = 95;
			9216: Pixel = 80;
			9217: Pixel = 70;
			9218: Pixel = 61;
			9219: Pixel = 62;
			9220: Pixel = 55;
			9221: Pixel = 52;
			9222: Pixel = 52;
			9223: Pixel = 82;
			9224: Pixel = 121;
			9225: Pixel = 129;
			9226: Pixel = 92;
			9227: Pixel = 68;
			9228: Pixel = 117;
			9229: Pixel = 130;
			9230: Pixel = 133;
			9231: Pixel = 139;
			9232: Pixel = 139;
			9233: Pixel = 136;
			9234: Pixel = 136;
			9235: Pixel = 138;
			9236: Pixel = 141;
			9237: Pixel = 143;
			9238: Pixel = 148;
			9239: Pixel = 153;
			9240: Pixel = 158;
			9241: Pixel = 162;
			9242: Pixel = 168;
			9243: Pixel = 175;
			9244: Pixel = 184;
			9245: Pixel = 191;
			9246: Pixel = 198;
			9247: Pixel = 204;
			9248: Pixel = 208;
			9249: Pixel = 211;
			9250: Pixel = 212;
			9251: Pixel = 231;
			9252: Pixel = 101;
			9253: Pixel = 55;
			9254: Pixel = 148;
			9255: Pixel = 148;
			9256: Pixel = 144;
			9257: Pixel = 143;
			9258: Pixel = 140;
			9259: Pixel = 139;
			9260: Pixel = 139;
			9261: Pixel = 136;
			9262: Pixel = 132;
			9263: Pixel = 126;
			9264: Pixel = 119;
			9265: Pixel = 168;
			9266: Pixel = 217;
			9267: Pixel = 206;
			9268: Pixel = 211;
			9269: Pixel = 218;
			9270: Pixel = 203;
			9271: Pixel = 142;
			9272: Pixel = 108;
			9273: Pixel = 99;
			9274: Pixel = 98;
			9275: Pixel = 112;
			9276: Pixel = 105;
			9277: Pixel = 90;
			9278: Pixel = 101;
			9279: Pixel = 103;
			9280: Pixel = 94;
			9281: Pixel = 83;
			9282: Pixel = 28;
			9283: Pixel = 52;
			9284: Pixel = 143;
			9285: Pixel = 176;
			9286: Pixel = 144;
			9287: Pixel = 48;
			9288: Pixel = 95;
			9289: Pixel = 165;
			9290: Pixel = 176;
			9291: Pixel = 175;
			9292: Pixel = 176;
			9293: Pixel = 166;
			9294: Pixel = 148;
			9295: Pixel = 92;
			9296: Pixel = 44;
			9297: Pixel = 47;
			9298: Pixel = 47;
			9299: Pixel = 48;
			9300: Pixel = 56;
			9301: Pixel = 47;
			9302: Pixel = 73;
			9303: Pixel = 64;
			9304: Pixel = 51;
			9305: Pixel = 55;
			9306: Pixel = 50;
			9307: Pixel = 46;
			9308: Pixel = 56;
			9309: Pixel = 78;
			9310: Pixel = 45;
			9311: Pixel = 65;
			9312: Pixel = 124;
			9313: Pixel = 122;
			9314: Pixel = 114;
			9315: Pixel = 54;
			9316: Pixel = 64;
			9317: Pixel = 75;
			9318: Pixel = 83;
			9319: Pixel = 95;
			9320: Pixel = 102;
			9321: Pixel = 82;
			9322: Pixel = 54;
			9323: Pixel = 49;
			9324: Pixel = 62;
			9325: Pixel = 97;
			9326: Pixel = 123;
			9327: Pixel = 132;
			9328: Pixel = 89;
			9329: Pixel = 77;
			9330: Pixel = 124;
			9331: Pixel = 132;
			9332: Pixel = 134;
			9333: Pixel = 139;
			9334: Pixel = 139;
			9335: Pixel = 137;
			9336: Pixel = 133;
			9337: Pixel = 135;
			9338: Pixel = 139;
			9339: Pixel = 142;
			9340: Pixel = 147;
			9341: Pixel = 151;
			9342: Pixel = 156;
			9343: Pixel = 159;
			9344: Pixel = 166;
			9345: Pixel = 171;
			9346: Pixel = 181;
			9347: Pixel = 189;
			9348: Pixel = 196;
			9349: Pixel = 202;
			9350: Pixel = 206;
			9351: Pixel = 210;
			9352: Pixel = 211;
			9353: Pixel = 228;
			9354: Pixel = 149;
			9355: Pixel = 69;
			9356: Pixel = 149;
			9357: Pixel = 147;
			9358: Pixel = 145;
			9359: Pixel = 142;
			9360: Pixel = 140;
			9361: Pixel = 138;
			9362: Pixel = 139;
			9363: Pixel = 137;
			9364: Pixel = 132;
			9365: Pixel = 126;
			9366: Pixel = 124;
			9367: Pixel = 176;
			9368: Pixel = 217;
			9369: Pixel = 203;
			9370: Pixel = 212;
			9371: Pixel = 217;
			9372: Pixel = 179;
			9373: Pixel = 121;
			9374: Pixel = 112;
			9375: Pixel = 98;
			9376: Pixel = 99;
			9377: Pixel = 108;
			9378: Pixel = 92;
			9379: Pixel = 91;
			9380: Pixel = 105;
			9381: Pixel = 98;
			9382: Pixel = 90;
			9383: Pixel = 90;
			9384: Pixel = 33;
			9385: Pixel = 45;
			9386: Pixel = 132;
			9387: Pixel = 175;
			9388: Pixel = 146;
			9389: Pixel = 55;
			9390: Pixel = 95;
			9391: Pixel = 162;
			9392: Pixel = 176;
			9393: Pixel = 177;
			9394: Pixel = 179;
			9395: Pixel = 167;
			9396: Pixel = 152;
			9397: Pixel = 87;
			9398: Pixel = 47;
			9399: Pixel = 46;
			9400: Pixel = 43;
			9401: Pixel = 55;
			9402: Pixel = 63;
			9403: Pixel = 49;
			9404: Pixel = 60;
			9405: Pixel = 59;
			9406: Pixel = 48;
			9407: Pixel = 55;
			9408: Pixel = 53;
			9409: Pixel = 44;
			9410: Pixel = 57;
			9411: Pixel = 79;
			9412: Pixel = 67;
			9413: Pixel = 91;
			9414: Pixel = 110;
			9415: Pixel = 110;
			9416: Pixel = 110;
			9417: Pixel = 112;
			9418: Pixel = 63;
			9419: Pixel = 40;
			9420: Pixel = 49;
			9421: Pixel = 53;
			9422: Pixel = 59;
			9423: Pixel = 68;
			9424: Pixel = 53;
			9425: Pixel = 47;
			9426: Pixel = 77;
			9427: Pixel = 107;
			9428: Pixel = 125;
			9429: Pixel = 130;
			9430: Pixel = 77;
			9431: Pixel = 90;
			9432: Pixel = 130;
			9433: Pixel = 135;
			9434: Pixel = 139;
			9435: Pixel = 139;
			9436: Pixel = 141;
			9437: Pixel = 139;
			9438: Pixel = 135;
			9439: Pixel = 136;
			9440: Pixel = 138;
			9441: Pixel = 140;
			9442: Pixel = 145;
			9443: Pixel = 149;
			9444: Pixel = 155;
			9445: Pixel = 158;
			9446: Pixel = 165;
			9447: Pixel = 169;
			9448: Pixel = 177;
			9449: Pixel = 187;
			9450: Pixel = 194;
			9451: Pixel = 200;
			9452: Pixel = 205;
			9453: Pixel = 208;
			9454: Pixel = 211;
			9455: Pixel = 220;
			9456: Pixel = 188;
			9457: Pixel = 94;
			9458: Pixel = 147;
			9459: Pixel = 148;
			9460: Pixel = 145;
			9461: Pixel = 143;
			9462: Pixel = 142;
			9463: Pixel = 140;
			9464: Pixel = 140;
			9465: Pixel = 137;
			9466: Pixel = 131;
			9467: Pixel = 130;
			9468: Pixel = 129;
			9469: Pixel = 157;
			9470: Pixel = 199;
			9471: Pixel = 199;
			9472: Pixel = 214;
			9473: Pixel = 213;
			9474: Pixel = 159;
			9475: Pixel = 112;
			9476: Pixel = 110;
			9477: Pixel = 96;
			9478: Pixel = 99;
			9479: Pixel = 90;
			9480: Pixel = 85;
			9481: Pixel = 103;
			9482: Pixel = 99;
			9483: Pixel = 93;
			9484: Pixel = 93;
			9485: Pixel = 95;
			9486: Pixel = 38;
			9487: Pixel = 39;
			9488: Pixel = 121;
			9489: Pixel = 172;
			9490: Pixel = 150;
			9491: Pixel = 70;
			9492: Pixel = 93;
			9493: Pixel = 161;
			9494: Pixel = 176;
			9495: Pixel = 175;
			9496: Pixel = 178;
			9497: Pixel = 165;
			9498: Pixel = 154;
			9499: Pixel = 107;
			9500: Pixel = 55;
			9501: Pixel = 40;
			9502: Pixel = 59;
			9503: Pixel = 70;
			9504: Pixel = 50;
			9505: Pixel = 45;
			9506: Pixel = 64;
			9507: Pixel = 54;
			9508: Pixel = 59;
			9509: Pixel = 56;
			9510: Pixel = 58;
			9511: Pixel = 51;
			9512: Pixel = 71;
			9513: Pixel = 59;
			9514: Pixel = 76;
			9515: Pixel = 71;
			9516: Pixel = 110;
			9517: Pixel = 119;
			9518: Pixel = 64;
			9519: Pixel = 109;
			9520: Pixel = 138;
			9521: Pixel = 74;
			9522: Pixel = 47;
			9523: Pixel = 55;
			9524: Pixel = 54;
			9525: Pixel = 47;
			9526: Pixel = 45;
			9527: Pixel = 55;
			9528: Pixel = 90;
			9529: Pixel = 115;
			9530: Pixel = 126;
			9531: Pixel = 117;
			9532: Pixel = 67;
			9533: Pixel = 105;
			9534: Pixel = 134;
			9535: Pixel = 138;
			9536: Pixel = 140;
			9537: Pixel = 143;
			9538: Pixel = 140;
			9539: Pixel = 138;
			9540: Pixel = 137;
			9541: Pixel = 135;
			9542: Pixel = 137;
			9543: Pixel = 141;
			9544: Pixel = 144;
			9545: Pixel = 148;
			9546: Pixel = 152;
			9547: Pixel = 156;
			9548: Pixel = 160;
			9549: Pixel = 166;
			9550: Pixel = 174;
			9551: Pixel = 183;
			9552: Pixel = 192;
			9553: Pixel = 198;
			9554: Pixel = 203;
			9555: Pixel = 208;
			9556: Pixel = 211;
			9557: Pixel = 213;
			9558: Pixel = 212;
			9559: Pixel = 142;
			9560: Pixel = 132;
			9561: Pixel = 126;
			9562: Pixel = 136;
			9563: Pixel = 141;
			9564: Pixel = 146;
			9565: Pixel = 145;
			9566: Pixel = 143;
			9567: Pixel = 140;
			9568: Pixel = 134;
			9569: Pixel = 136;
			9570: Pixel = 141;
			9571: Pixel = 139;
			9572: Pixel = 144;
			9573: Pixel = 187;
			9574: Pixel = 220;
			9575: Pixel = 206;
			9576: Pixel = 144;
			9577: Pixel = 108;
			9578: Pixel = 99;
			9579: Pixel = 93;
			9580: Pixel = 97;
			9581: Pixel = 77;
			9582: Pixel = 97;
			9583: Pixel = 105;
			9584: Pixel = 89;
			9585: Pixel = 90;
			9586: Pixel = 97;
			9587: Pixel = 89;
			9588: Pixel = 36;
			9589: Pixel = 38;
			9590: Pixel = 116;
			9591: Pixel = 169;
			9592: Pixel = 153;
			9593: Pixel = 75;
			9594: Pixel = 91;
			9595: Pixel = 158;
			9596: Pixel = 174;
			9597: Pixel = 175;
			9598: Pixel = 178;
			9599: Pixel = 168;
			9600: Pixel = 145;
			9601: Pixel = 104;
			9602: Pixel = 59;
			9603: Pixel = 43;
			9604: Pixel = 54;
			9605: Pixel = 48;
			9606: Pixel = 45;
			9607: Pixel = 56;
			9608: Pixel = 60;
			9609: Pixel = 61;
			9610: Pixel = 63;
			9611: Pixel = 49;
			9612: Pixel = 51;
			9613: Pixel = 48;
			9614: Pixel = 65;
			9615: Pixel = 49;
			9616: Pixel = 107;
			9617: Pixel = 72;
			9618: Pixel = 39;
			9619: Pixel = 87;
			9620: Pixel = 69;
			9621: Pixel = 85;
			9622: Pixel = 129;
			9623: Pixel = 56;
			9624: Pixel = 46;
			9625: Pixel = 50;
			9626: Pixel = 49;
			9627: Pixel = 43;
			9628: Pixel = 48;
			9629: Pixel = 67;
			9630: Pixel = 102;
			9631: Pixel = 118;
			9632: Pixel = 129;
			9633: Pixel = 95;
			9634: Pixel = 67;
			9635: Pixel = 125;
			9636: Pixel = 136;
			9637: Pixel = 137;
			9638: Pixel = 140;
			9639: Pixel = 143;
			9640: Pixel = 142;
			9641: Pixel = 141;
			9642: Pixel = 140;
			9643: Pixel = 136;
			9644: Pixel = 138;
			9645: Pixel = 140;
			9646: Pixel = 144;
			9647: Pixel = 148;
			9648: Pixel = 151;
			9649: Pixel = 153;
			9650: Pixel = 159;
			9651: Pixel = 164;
			9652: Pixel = 171;
			9653: Pixel = 179;
			9654: Pixel = 189;
			9655: Pixel = 195;
			9656: Pixel = 202;
			9657: Pixel = 208;
			9658: Pixel = 211;
			9659: Pixel = 211;
			9660: Pixel = 220;
			9661: Pixel = 175;
			9662: Pixel = 94;
			9663: Pixel = 85;
			9664: Pixel = 97;
			9665: Pixel = 112;
			9666: Pixel = 125;
			9667: Pixel = 135;
			9668: Pixel = 140;
			9669: Pixel = 141;
			9670: Pixel = 140;
			9671: Pixel = 147;
			9672: Pixel = 151;
			9673: Pixel = 136;
			9674: Pixel = 136;
			9675: Pixel = 195;
			9676: Pixel = 222;
			9677: Pixel = 192;
			9678: Pixel = 127;
			9679: Pixel = 100;
			9680: Pixel = 88;
			9681: Pixel = 98;
			9682: Pixel = 79;
			9683: Pixel = 86;
			9684: Pixel = 103;
			9685: Pixel = 95;
			9686: Pixel = 90;
			9687: Pixel = 98;
			9688: Pixel = 92;
			9689: Pixel = 70;
			9690: Pixel = 34;
			9691: Pixel = 32;
			9692: Pixel = 106;
			9693: Pixel = 177;
			9694: Pixel = 165;
			9695: Pixel = 82;
			9696: Pixel = 86;
			9697: Pixel = 155;
			9698: Pixel = 172;
			9699: Pixel = 175;
			9700: Pixel = 178;
			9701: Pixel = 171;
			9702: Pixel = 142;
			9703: Pixel = 101;
			9704: Pixel = 67;
			9705: Pixel = 44;
			9706: Pixel = 51;
			9707: Pixel = 43;
			9708: Pixel = 54;
			9709: Pixel = 60;
			9710: Pixel = 55;
			9711: Pixel = 58;
			9712: Pixel = 65;
			9713: Pixel = 45;
			9714: Pixel = 44;
			9715: Pixel = 48;
			9716: Pixel = 54;
			9717: Pixel = 74;
			9718: Pixel = 114;
			9719: Pixel = 117;
			9720: Pixel = 61;
			9721: Pixel = 59;
			9722: Pixel = 75;
			9723: Pixel = 91;
			9724: Pixel = 71;
			9725: Pixel = 46;
			9726: Pixel = 45;
			9727: Pixel = 47;
			9728: Pixel = 44;
			9729: Pixel = 41;
			9730: Pixel = 59;
			9731: Pixel = 86;
			9732: Pixel = 115;
			9733: Pixel = 118;
			9734: Pixel = 121;
			9735: Pixel = 61;
			9736: Pixel = 89;
			9737: Pixel = 134;
			9738: Pixel = 134;
			9739: Pixel = 137;
			9740: Pixel = 142;
			9741: Pixel = 143;
			9742: Pixel = 140;
			9743: Pixel = 141;
			9744: Pixel = 139;
			9745: Pixel = 137;
			9746: Pixel = 135;
			9747: Pixel = 137;
			9748: Pixel = 142;
			9749: Pixel = 145;
			9750: Pixel = 149;
			9751: Pixel = 153;
			9752: Pixel = 158;
			9753: Pixel = 163;
			9754: Pixel = 169;
			9755: Pixel = 174;
			9756: Pixel = 186;
			9757: Pixel = 192;
			9758: Pixel = 201;
			9759: Pixel = 207;
			9760: Pixel = 211;
			9761: Pixel = 211;
			9762: Pixel = 222;
			9763: Pixel = 188;
			9764: Pixel = 75;
			9765: Pixel = 79;
			9766: Pixel = 74;
			9767: Pixel = 79;
			9768: Pixel = 84;
			9769: Pixel = 91;
			9770: Pixel = 101;
			9771: Pixel = 110;
			9772: Pixel = 129;
			9773: Pixel = 153;
			9774: Pixel = 151;
			9775: Pixel = 134;
			9776: Pixel = 152;
			9777: Pixel = 212;
			9778: Pixel = 216;
			9779: Pixel = 164;
			9780: Pixel = 104;
			9781: Pixel = 76;
			9782: Pixel = 86;
			9783: Pixel = 88;
			9784: Pixel = 77;
			9785: Pixel = 101;
			9786: Pixel = 96;
			9787: Pixel = 91;
			9788: Pixel = 97;
			9789: Pixel = 102;
			9790: Pixel = 82;
			9791: Pixel = 57;
			9792: Pixel = 38;
			9793: Pixel = 32;
			9794: Pixel = 103;
			9795: Pixel = 177;
			9796: Pixel = 173;
			9797: Pixel = 97;
			9798: Pixel = 83;
			9799: Pixel = 154;
			9800: Pixel = 172;
			9801: Pixel = 175;
			9802: Pixel = 178;
			9803: Pixel = 176;
			9804: Pixel = 129;
			9805: Pixel = 98;
			9806: Pixel = 66;
			9807: Pixel = 45;
			9808: Pixel = 42;
			9809: Pixel = 48;
			9810: Pixel = 61;
			9811: Pixel = 52;
			9812: Pixel = 54;
			9813: Pixel = 57;
			9814: Pixel = 64;
			9815: Pixel = 57;
			9816: Pixel = 48;
			9817: Pixel = 51;
			9818: Pixel = 52;
			9819: Pixel = 44;
			9820: Pixel = 80;
			9821: Pixel = 136;
			9822: Pixel = 118;
			9823: Pixel = 94;
			9824: Pixel = 99;
			9825: Pixel = 50;
			9826: Pixel = 45;
			9827: Pixel = 51;
			9828: Pixel = 46;
			9829: Pixel = 43;
			9830: Pixel = 40;
			9831: Pixel = 45;
			9832: Pixel = 71;
			9833: Pixel = 102;
			9834: Pixel = 116;
			9835: Pixel = 125;
			9836: Pixel = 79;
			9837: Pixel = 54;
			9838: Pixel = 121;
			9839: Pixel = 136;
			9840: Pixel = 135;
			9841: Pixel = 138;
			9842: Pixel = 139;
			9843: Pixel = 140;
			9844: Pixel = 142;
			9845: Pixel = 142;
			9846: Pixel = 139;
			9847: Pixel = 138;
			9848: Pixel = 135;
			9849: Pixel = 136;
			9850: Pixel = 139;
			9851: Pixel = 143;
			9852: Pixel = 147;
			9853: Pixel = 151;
			9854: Pixel = 155;
			9855: Pixel = 160;
			9856: Pixel = 165;
			9857: Pixel = 172;
			9858: Pixel = 182;
			9859: Pixel = 190;
			9860: Pixel = 198;
			9861: Pixel = 204;
			9862: Pixel = 209;
			9863: Pixel = 211;
			9864: Pixel = 217;
			9865: Pixel = 210;
			9866: Pixel = 96;
			9867: Pixel = 93;
			9868: Pixel = 94;
			9869: Pixel = 86;
			9870: Pixel = 75;
			9871: Pixel = 64;
			9872: Pixel = 58;
			9873: Pixel = 54;
			9874: Pixel = 71;
			9875: Pixel = 109;
			9876: Pixel = 167;
			9877: Pixel = 172;
			9878: Pixel = 170;
			9879: Pixel = 217;
			9880: Pixel = 202;
			9881: Pixel = 127;
			9882: Pixel = 68;
			9883: Pixel = 67;
			9884: Pixel = 83;
			9885: Pixel = 78;
			9886: Pixel = 100;
			9887: Pixel = 99;
			9888: Pixel = 88;
			9889: Pixel = 91;
			9890: Pixel = 100;
			9891: Pixel = 97;
			9892: Pixel = 70;
			9893: Pixel = 52;
			9894: Pixel = 71;
			9895: Pixel = 69;
			9896: Pixel = 105;
			9897: Pixel = 175;
			9898: Pixel = 182;
			9899: Pixel = 107;
			9900: Pixel = 86;
			9901: Pixel = 153;
			9902: Pixel = 173;
			9903: Pixel = 174;
			9904: Pixel = 179;
			9905: Pixel = 176;
			9906: Pixel = 125;
			9907: Pixel = 102;
			9908: Pixel = 51;
			9909: Pixel = 47;
			9910: Pixel = 55;
			9911: Pixel = 52;
			9912: Pixel = 51;
			9913: Pixel = 50;
			9914: Pixel = 54;
			9915: Pixel = 61;
			9916: Pixel = 61;
			9917: Pixel = 57;
			9918: Pixel = 49;
			9919: Pixel = 43;
			9920: Pixel = 51;
			9921: Pixel = 57;
			9922: Pixel = 44;
			9923: Pixel = 89;
			9924: Pixel = 146;
			9925: Pixel = 113;
			9926: Pixel = 102;
			9927: Pixel = 73;
			9928: Pixel = 43;
			9929: Pixel = 45;
			9930: Pixel = 44;
			9931: Pixel = 41;
			9932: Pixel = 40;
			9933: Pixel = 57;
			9934: Pixel = 87;
			9935: Pixel = 111;
			9936: Pixel = 124;
			9937: Pixel = 101;
			9938: Pixel = 42;
			9939: Pixel = 97;
			9940: Pixel = 134;
			9941: Pixel = 134;
			9942: Pixel = 137;
			9943: Pixel = 138;
			9944: Pixel = 139;
			9945: Pixel = 140;
			9946: Pixel = 143;
			9947: Pixel = 143;
			9948: Pixel = 142;
			9949: Pixel = 139;
			9950: Pixel = 137;
			9951: Pixel = 137;
			9952: Pixel = 138;
			9953: Pixel = 139;
			9954: Pixel = 144;
			9955: Pixel = 148;
			9956: Pixel = 154;
			9957: Pixel = 156;
			9958: Pixel = 161;
			9959: Pixel = 171;
			9960: Pixel = 178;
			9961: Pixel = 187;
			9962: Pixel = 196;
			9963: Pixel = 202;
			9964: Pixel = 207;
			9965: Pixel = 210;
			9966: Pixel = 212;
			9967: Pixel = 223;
			9968: Pixel = 129;
			9969: Pixel = 90;
			9970: Pixel = 108;
			9971: Pixel = 101;
			9972: Pixel = 91;
			9973: Pixel = 79;
			9974: Pixel = 60;
			9975: Pixel = 45;
			9976: Pixel = 29;
			9977: Pixel = 96;
			9978: Pixel = 208;
			9979: Pixel = 171;
			9980: Pixel = 183;
			9981: Pixel = 221;
			9982: Pixel = 170;
			9983: Pixel = 75;
			9984: Pixel = 59;
			9985: Pixel = 77;
			9986: Pixel = 72;
			9987: Pixel = 91;
			9988: Pixel = 106;
			9989: Pixel = 87;
			9990: Pixel = 82;
			9991: Pixel = 92;
			9992: Pixel = 108;
			9993: Pixel = 89;
			9994: Pixel = 65;
			9995: Pixel = 54;
			9996: Pixel = 92;
			9997: Pixel = 92;
			9998: Pixel = 120;
			9999: Pixel = 171;
			10000: Pixel = 185;
			10001: Pixel = 123;
			10002: Pixel = 90;
			10003: Pixel = 150;
			10004: Pixel = 174;
			10005: Pixel = 176;
			10006: Pixel = 181;
			10007: Pixel = 175;
			10008: Pixel = 123;
			10009: Pixel = 103;
			10010: Pixel = 51;
			10011: Pixel = 47;
			10012: Pixel = 52;
			10013: Pixel = 46;
			10014: Pixel = 50;
			10015: Pixel = 52;
			10016: Pixel = 49;
			10017: Pixel = 54;
			10018: Pixel = 62;
			10019: Pixel = 59;
			10020: Pixel = 48;
			10021: Pixel = 47;
			10022: Pixel = 52;
			10023: Pixel = 62;
			10024: Pixel = 54;
			10025: Pixel = 58;
			10026: Pixel = 93;
			10027: Pixel = 123;
			10028: Pixel = 110;
			10029: Pixel = 63;
			10030: Pixel = 44;
			10031: Pixel = 45;
			10032: Pixel = 41;
			10033: Pixel = 38;
			10034: Pixel = 49;
			10035: Pixel = 74;
			10036: Pixel = 104;
			10037: Pixel = 126;
			10038: Pixel = 99;
			10039: Pixel = 43;
			10040: Pixel = 81;
			10041: Pixel = 127;
			10042: Pixel = 131;
			10043: Pixel = 134;
			10044: Pixel = 138;
			10045: Pixel = 139;
			10046: Pixel = 138;
			10047: Pixel = 139;
			10048: Pixel = 142;
			10049: Pixel = 142;
			10050: Pixel = 142;
			10051: Pixel = 140;
			10052: Pixel = 139;
			10053: Pixel = 136;
			10054: Pixel = 139;
			10055: Pixel = 139;
			10056: Pixel = 142;
			10057: Pixel = 146;
			10058: Pixel = 151;
			10059: Pixel = 154;
			10060: Pixel = 161;
			10061: Pixel = 165;
			10062: Pixel = 173;
			10063: Pixel = 184;
			10064: Pixel = 193;
			10065: Pixel = 199;
			10066: Pixel = 206;
			10067: Pixel = 209;
			10068: Pixel = 210;
			10069: Pixel = 223;
			10070: Pixel = 164;
			10071: Pixel = 82;
			10072: Pixel = 109;
			10073: Pixel = 107;
			10074: Pixel = 98;
			10075: Pixel = 90;
			10076: Pixel = 79;
			10077: Pixel = 62;
			10078: Pixel = 39;
			10079: Pixel = 100;
			10080: Pixel = 201;
			10081: Pixel = 184;
			10082: Pixel = 196;
			10083: Pixel = 185;
			10084: Pixel = 88;
			10085: Pixel = 48;
			10086: Pixel = 69;
			10087: Pixel = 69;
			10088: Pixel = 82;
			10089: Pixel = 106;
			10090: Pixel = 88;
			10091: Pixel = 75;
			10092: Pixel = 82;
			10093: Pixel = 105;
			10094: Pixel = 107;
			10095: Pixel = 87;
			10096: Pixel = 70;
			10097: Pixel = 61;
			10098: Pixel = 83;
			10099: Pixel = 108;
			10100: Pixel = 128;
			10101: Pixel = 169;
			10102: Pixel = 181;
			10103: Pixel = 129;
			10104: Pixel = 93;
			10105: Pixel = 149;
			10106: Pixel = 173;
			10107: Pixel = 176;
			10108: Pixel = 182;
			10109: Pixel = 176;
			10110: Pixel = 120;
			10111: Pixel = 96;
			10112: Pixel = 46;
			10113: Pixel = 49;
			10114: Pixel = 49;
			10115: Pixel = 51;
			10116: Pixel = 52;
			10117: Pixel = 54;
			10118: Pixel = 43;
			10119: Pixel = 65;
			10120: Pixel = 64;
			10121: Pixel = 68;
			10122: Pixel = 64;
			10123: Pixel = 42;
			10124: Pixel = 75;
			10125: Pixel = 61;
			10126: Pixel = 65;
			10127: Pixel = 68;
			10128: Pixel = 87;
			10129: Pixel = 98;
			10130: Pixel = 81;
			10131: Pixel = 52;
			10132: Pixel = 44;
			10133: Pixel = 45;
			10134: Pixel = 38;
			10135: Pixel = 43;
			10136: Pixel = 70;
			10137: Pixel = 94;
			10138: Pixel = 100;
			10139: Pixel = 74;
			10140: Pixel = 48;
			10141: Pixel = 82;
			10142: Pixel = 119;
			10143: Pixel = 127;
			10144: Pixel = 131;
			10145: Pixel = 135;
			10146: Pixel = 138;
			10147: Pixel = 138;
			10148: Pixel = 139;
			10149: Pixel = 139;
			10150: Pixel = 142;
			10151: Pixel = 142;
			10152: Pixel = 143;
			10153: Pixel = 143;
			10154: Pixel = 141;
			10155: Pixel = 139;
			10156: Pixel = 140;
			10157: Pixel = 138;
			10158: Pixel = 140;
			10159: Pixel = 145;
			10160: Pixel = 147;
			10161: Pixel = 152;
			10162: Pixel = 159;
			10163: Pixel = 164;
			10164: Pixel = 169;
			10165: Pixel = 176;
			10166: Pixel = 187;
			10167: Pixel = 195;
			10168: Pixel = 203;
			10169: Pixel = 208;
			10170: Pixel = 210;
			10171: Pixel = 217;
			10172: Pixel = 196;
			10173: Pixel = 87;
			10174: Pixel = 99;
			10175: Pixel = 106;
			10176: Pixel = 100;
			10177: Pixel = 96;
			10178: Pixel = 89;
			10179: Pixel = 80;
			10180: Pixel = 74;
			10181: Pixel = 107;
			10182: Pixel = 201;
			10183: Pixel = 209;
			10184: Pixel = 154;
			10185: Pixel = 90;
			10186: Pixel = 53;
			10187: Pixel = 66;
			10188: Pixel = 68;
			10189: Pixel = 77;
			10190: Pixel = 105;
			10191: Pixel = 96;
			10192: Pixel = 74;
			10193: Pixel = 76;
			10194: Pixel = 96;
			10195: Pixel = 112;
			10196: Pixel = 98;
			10197: Pixel = 81;
			10198: Pixel = 64;
			10199: Pixel = 67;
			10200: Pixel = 65;
			10201: Pixel = 98;
			10202: Pixel = 110;
			10203: Pixel = 160;
			10204: Pixel = 180;
			10205: Pixel = 133;
			10206: Pixel = 95;
			10207: Pixel = 146;
			10208: Pixel = 173;
			10209: Pixel = 178;
			10210: Pixel = 181;
			10211: Pixel = 178;
			10212: Pixel = 122;
			10213: Pixel = 77;
			10214: Pixel = 42;
			10215: Pixel = 50;
			10216: Pixel = 53;
			10217: Pixel = 56;
			10218: Pixel = 51;
			10219: Pixel = 61;
			10220: Pixel = 44;
			10221: Pixel = 72;
			10222: Pixel = 71;
			10223: Pixel = 72;
			10224: Pixel = 94;
			10225: Pixel = 48;
			10226: Pixel = 69;
			10227: Pixel = 52;
			10228: Pixel = 84;
			10229: Pixel = 62;
			10230: Pixel = 86;
			10231: Pixel = 131;
			10232: Pixel = 69;
			10233: Pixel = 50;
			10234: Pixel = 41;
			10235: Pixel = 45;
			10236: Pixel = 43;
			10237: Pixel = 46;
			10238: Pixel = 60;
			10239: Pixel = 59;
			10240: Pixel = 56;
			10241: Pixel = 69;
			10242: Pixel = 103;
			10243: Pixel = 122;
			10244: Pixel = 123;
			10245: Pixel = 128;
			10246: Pixel = 131;
			10247: Pixel = 135;
			10248: Pixel = 136;
			10249: Pixel = 138;
			10250: Pixel = 139;
			10251: Pixel = 139;
			10252: Pixel = 141;
			10253: Pixel = 143;
			10254: Pixel = 145;
			10255: Pixel = 146;
			10256: Pixel = 143;
			10257: Pixel = 142;
			10258: Pixel = 139;
			10259: Pixel = 140;
			10260: Pixel = 140;
			10261: Pixel = 143;
			10262: Pixel = 147;
			10263: Pixel = 151;
			10264: Pixel = 156;
			10265: Pixel = 162;
			10266: Pixel = 169;
			10267: Pixel = 176;
			10268: Pixel = 183;
			10269: Pixel = 192;
			10270: Pixel = 200;
			10271: Pixel = 206;
			10272: Pixel = 210;
			10273: Pixel = 213;
			10274: Pixel = 215;
			10275: Pixel = 107;
			10276: Pixel = 87;
			10277: Pixel = 102;
			10278: Pixel = 103;
			10279: Pixel = 102;
			10280: Pixel = 97;
			10281: Pixel = 98;
			10282: Pixel = 99;
			10283: Pixel = 110;
			10284: Pixel = 181;
			10285: Pixel = 156;
			10286: Pixel = 83;
			10287: Pixel = 68;
			10288: Pixel = 73;
			10289: Pixel = 75;
			10290: Pixel = 77;
			10291: Pixel = 106;
			10292: Pixel = 101;
			10293: Pixel = 77;
			10294: Pixel = 65;
			10295: Pixel = 84;
			10296: Pixel = 110;
			10297: Pixel = 110;
			10298: Pixel = 95;
			10299: Pixel = 68;
			10300: Pixel = 66;
			10301: Pixel = 62;
			10302: Pixel = 52;
			10303: Pixel = 73;
			10304: Pixel = 97;
			10305: Pixel = 152;
			10306: Pixel = 178;
			10307: Pixel = 139;
			10308: Pixel = 101;
			10309: Pixel = 143;
			10310: Pixel = 173;
			10311: Pixel = 179;
			10312: Pixel = 181;
			10313: Pixel = 180;
			10314: Pixel = 125;
			10315: Pixel = 55;
			10316: Pixel = 47;
			10317: Pixel = 49;
			10318: Pixel = 51;
			10319: Pixel = 61;
			10320: Pixel = 57;
			10321: Pixel = 68;
			10322: Pixel = 45;
			10323: Pixel = 70;
			10324: Pixel = 60;
			10325: Pixel = 65;
			10326: Pixel = 117;
			10327: Pixel = 57;
			10328: Pixel = 71;
			10329: Pixel = 73;
			10330: Pixel = 58;
			10331: Pixel = 83;
			10332: Pixel = 80;
			10333: Pixel = 119;
			10334: Pixel = 96;
			10335: Pixel = 49;
			10336: Pixel = 46;
			10337: Pixel = 44;
			10338: Pixel = 43;
			10339: Pixel = 50;
			10340: Pixel = 64;
			10341: Pixel = 81;
			10342: Pixel = 100;
			10343: Pixel = 118;
			10344: Pixel = 122;
			10345: Pixel = 124;
			10346: Pixel = 128;
			10347: Pixel = 127;
			10348: Pixel = 128;
			10349: Pixel = 132;
			10350: Pixel = 135;
			10351: Pixel = 136;
			10352: Pixel = 137;
			10353: Pixel = 141;
			10354: Pixel = 141;
			10355: Pixel = 142;
			10356: Pixel = 145;
			10357: Pixel = 145;
			10358: Pixel = 143;
			10359: Pixel = 144;
			10360: Pixel = 142;
			10361: Pixel = 141;
			10362: Pixel = 142;
			10363: Pixel = 142;
			10364: Pixel = 146;
			10365: Pixel = 150;
			10366: Pixel = 155;
			10367: Pixel = 159;
			10368: Pixel = 166;
			10369: Pixel = 174;
			10370: Pixel = 182;
			10371: Pixel = 188;
			10372: Pixel = 195;
			10373: Pixel = 202;
			10374: Pixel = 209;
			10375: Pixel = 210;
			10376: Pixel = 223;
			10377: Pixel = 137;
			10378: Pixel = 75;
			10379: Pixel = 98;
			10380: Pixel = 104;
			10381: Pixel = 109;
			10382: Pixel = 104;
			10383: Pixel = 113;
			10384: Pixel = 114;
			10385: Pixel = 110;
			10386: Pixel = 114;
			10387: Pixel = 93;
			10388: Pixel = 84;
			10389: Pixel = 92;
			10390: Pixel = 84;
			10391: Pixel = 73;
			10392: Pixel = 95;
			10393: Pixel = 102;
			10394: Pixel = 81;
			10395: Pixel = 66;
			10396: Pixel = 70;
			10397: Pixel = 104;
			10398: Pixel = 117;
			10399: Pixel = 110;
			10400: Pixel = 85;
			10401: Pixel = 63;
			10402: Pixel = 60;
			10403: Pixel = 53;
			10404: Pixel = 56;
			10405: Pixel = 60;
			10406: Pixel = 77;
			10407: Pixel = 156;
			10408: Pixel = 199;
			10409: Pixel = 165;
			10410: Pixel = 108;
			10411: Pixel = 143;
			10412: Pixel = 174;
			10413: Pixel = 179;
			10414: Pixel = 184;
			10415: Pixel = 176;
			10416: Pixel = 95;
			10417: Pixel = 55;
			10418: Pixel = 52;
			10419: Pixel = 48;
			10420: Pixel = 51;
			10421: Pixel = 59;
			10422: Pixel = 55;
			10423: Pixel = 70;
			10424: Pixel = 47;
			10425: Pixel = 75;
			10426: Pixel = 57;
			10427: Pixel = 60;
			10428: Pixel = 103;
			10429: Pixel = 89;
			10430: Pixel = 56;
			10431: Pixel = 102;
			10432: Pixel = 39;
			10433: Pixel = 87;
			10434: Pixel = 69;
			10435: Pixel = 95;
			10436: Pixel = 83;
			10437: Pixel = 43;
			10438: Pixel = 44;
			10439: Pixel = 46;
			10440: Pixel = 51;
			10441: Pixel = 78;
			10442: Pixel = 101;
			10443: Pixel = 114;
			10444: Pixel = 115;
			10445: Pixel = 120;
			10446: Pixel = 125;
			10447: Pixel = 126;
			10448: Pixel = 128;
			10449: Pixel = 128;
			10450: Pixel = 129;
			10451: Pixel = 133;
			10452: Pixel = 135;
			10453: Pixel = 135;
			10454: Pixel = 138;
			10455: Pixel = 139;
			10456: Pixel = 140;
			10457: Pixel = 141;
			10458: Pixel = 143;
			10459: Pixel = 144;
			10460: Pixel = 146;
			10461: Pixel = 145;
			10462: Pixel = 146;
			10463: Pixel = 144;
			10464: Pixel = 143;
			10465: Pixel = 145;
			10466: Pixel = 147;
			10467: Pixel = 149;
			10468: Pixel = 152;
			10469: Pixel = 158;
			10470: Pixel = 165;
			10471: Pixel = 170;
			10472: Pixel = 178;
			10473: Pixel = 184;
			10474: Pixel = 191;
			10475: Pixel = 199;
			10476: Pixel = 206;
			10477: Pixel = 207;
			10478: Pixel = 219;
			10479: Pixel = 167;
			10480: Pixel = 72;
			10481: Pixel = 96;
			10482: Pixel = 105;
			10483: Pixel = 110;
			10484: Pixel = 117;
			10485: Pixel = 119;
			10486: Pixel = 115;
			10487: Pixel = 113;
			10488: Pixel = 103;
			10489: Pixel = 98;
			10490: Pixel = 109;
			10491: Pixel = 104;
			10492: Pixel = 84;
			10493: Pixel = 90;
			10494: Pixel = 97;
			10495: Pixel = 75;
			10496: Pixel = 72;
			10497: Pixel = 71;
			10498: Pixel = 90;
			10499: Pixel = 120;
			10500: Pixel = 117;
			10501: Pixel = 97;
			10502: Pixel = 70;
			10503: Pixel = 58;
			10504: Pixel = 54;
			10505: Pixel = 51;
			10506: Pixel = 52;
			10507: Pixel = 52;
			10508: Pixel = 69;
			10509: Pixel = 173;
			10510: Pixel = 208;
			10511: Pixel = 191;
			10512: Pixel = 121;
			10513: Pixel = 140;
			10514: Pixel = 174;
			10515: Pixel = 177;
			10516: Pixel = 182;
			10517: Pixel = 173;
			10518: Pixel = 107;
			10519: Pixel = 51;
			10520: Pixel = 51;
			10521: Pixel = 50;
			10522: Pixel = 57;
			10523: Pixel = 57;
			10524: Pixel = 66;
			10525: Pixel = 64;
			10526: Pixel = 55;
			10527: Pixel = 89;
			10528: Pixel = 59;
			10529: Pixel = 74;
			10530: Pixel = 86;
			10531: Pixel = 113;
			10532: Pixel = 54;
			10533: Pixel = 82;
			10534: Pixel = 62;
			10535: Pixel = 68;
			10536: Pixel = 76;
			10537: Pixel = 66;
			10538: Pixel = 100;
			10539: Pixel = 77;
			10540: Pixel = 34;
			10541: Pixel = 51;
			10542: Pixel = 75;
			10543: Pixel = 98;
			10544: Pixel = 109;
			10545: Pixel = 115;
			10546: Pixel = 118;
			10547: Pixel = 120;
			10548: Pixel = 126;
			10549: Pixel = 126;
			10550: Pixel = 127;
			10551: Pixel = 131;
			10552: Pixel = 131;
			10553: Pixel = 131;
			10554: Pixel = 134;
			10555: Pixel = 136;
			10556: Pixel = 136;
			10557: Pixel = 139;
			10558: Pixel = 139;
			10559: Pixel = 140;
			10560: Pixel = 143;
			10561: Pixel = 145;
			10562: Pixel = 146;
			10563: Pixel = 146;
			10564: Pixel = 147;
			10565: Pixel = 148;
			10566: Pixel = 147;
			10567: Pixel = 146;
			10568: Pixel = 148;
			10569: Pixel = 152;
			10570: Pixel = 152;
			10571: Pixel = 159;
			10572: Pixel = 165;
			10573: Pixel = 168;
			10574: Pixel = 176;
			10575: Pixel = 182;
			10576: Pixel = 189;
			10577: Pixel = 197;
			10578: Pixel = 203;
			10579: Pixel = 206;
			10580: Pixel = 214;
			10581: Pixel = 196;
			10582: Pixel = 81;
			10583: Pixel = 89;
			10584: Pixel = 100;
			10585: Pixel = 107;
			10586: Pixel = 118;
			10587: Pixel = 120;
			10588: Pixel = 119;
			10589: Pixel = 114;
			10590: Pixel = 112;
			10591: Pixel = 118;
			10592: Pixel = 122;
			10593: Pixel = 101;
			10594: Pixel = 94;
			10595: Pixel = 96;
			10596: Pixel = 85;
			10597: Pixel = 78;
			10598: Pixel = 74;
			10599: Pixel = 86;
			10600: Pixel = 118;
			10601: Pixel = 124;
			10602: Pixel = 105;
			10603: Pixel = 77;
			10604: Pixel = 54;
			10605: Pixel = 54;
			10606: Pixel = 59;
			10607: Pixel = 77;
			10608: Pixel = 49;
			10609: Pixel = 51;
			10610: Pixel = 60;
			10611: Pixel = 169;
			10612: Pixel = 203;
			10613: Pixel = 188;
			10614: Pixel = 123;
			10615: Pixel = 141;
			10616: Pixel = 173;
			10617: Pixel = 178;
			10618: Pixel = 182;
			10619: Pixel = 170;
			10620: Pixel = 92;
			10621: Pixel = 51;
			10622: Pixel = 45;
			10623: Pixel = 53;
			10624: Pixel = 57;
			10625: Pixel = 64;
			10626: Pixel = 73;
			10627: Pixel = 64;
			10628: Pixel = 71;
			10629: Pixel = 100;
			10630: Pixel = 51;
			10631: Pixel = 80;
			10632: Pixel = 74;
			10633: Pixel = 84;
			10634: Pixel = 87;
			10635: Pixel = 91;
			10636: Pixel = 68;
			10637: Pixel = 53;
			10638: Pixel = 73;
			10639: Pixel = 53;
			10640: Pixel = 76;
			10641: Pixel = 98;
			10642: Pixel = 71;
			10643: Pixel = 68;
			10644: Pixel = 88;
			10645: Pixel = 100;
			10646: Pixel = 111;
			10647: Pixel = 117;
			10648: Pixel = 121;
			10649: Pixel = 123;
			10650: Pixel = 126;
			10651: Pixel = 126;
			10652: Pixel = 128;
			10653: Pixel = 129;
			10654: Pixel = 131;
			10655: Pixel = 130;
			10656: Pixel = 135;
			10657: Pixel = 137;
			10658: Pixel = 133;
			10659: Pixel = 137;
			10660: Pixel = 139;
			10661: Pixel = 140;
			10662: Pixel = 144;
			10663: Pixel = 145;
			10664: Pixel = 143;
			10665: Pixel = 145;
			10666: Pixel = 146;
			10667: Pixel = 149;
			10668: Pixel = 148;
			10669: Pixel = 148;
			10670: Pixel = 149;
			10671: Pixel = 152;
			10672: Pixel = 156;
			10673: Pixel = 159;
			10674: Pixel = 164;
			10675: Pixel = 166;
			10676: Pixel = 172;
			10677: Pixel = 180;
			10678: Pixel = 188;
			10679: Pixel = 194;
			10680: Pixel = 200;
			10681: Pixel = 205;
			10682: Pixel = 209;
			10683: Pixel = 212;
			10684: Pixel = 115;
			10685: Pixel = 86;
			10686: Pixel = 93;
			10687: Pixel = 103;
			10688: Pixel = 113;
			10689: Pixel = 127;
			10690: Pixel = 126;
			10691: Pixel = 120;
			10692: Pixel = 127;
			10693: Pixel = 136;
			10694: Pixel = 118;
			10695: Pixel = 94;
			10696: Pixel = 86;
			10697: Pixel = 77;
			10698: Pixel = 85;
			10699: Pixel = 88;
			10700: Pixel = 82;
			10701: Pixel = 107;
			10702: Pixel = 130;
			10703: Pixel = 120;
			10704: Pixel = 83;
			10705: Pixel = 55;
			10706: Pixel = 46;
			10707: Pixel = 54;
			10708: Pixel = 80;
			10709: Pixel = 101;
		endcase
	end
endmodule